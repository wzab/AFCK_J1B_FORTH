
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;

package ram_prog is

type T_RAM_PROG is array(0 to 8191) of std_logic_vector(31 downto 0);
constant ram_init : T_RAM_PROG := (
  0 => std_logic_vector'(x"45f145fc"),
  1 => std_logic_vector'(x"628f8001"),
  2 => std_logic_vector'(x"66008000"),
  3 => std_logic_vector'(x"8000628f"),
  4 => std_logic_vector'(x"8004678f"),
  5 => std_logic_vector'(x"8002628f"),
  6 => std_logic_vector'(x"67036a8f"),
  7 => std_logic_vector'(x"6110668c"),
  8 => std_logic_vector'(x"8000688f"),
  9 => std_logic_vector'(x"8000688f"),
  10 => std_logic_vector'(x"8000000f"),
  11 => std_logic_vector'(x"6110000d"),
  12 => std_logic_vector'(x"80006f8f"),
  13 => std_logic_vector'(x"60336110"),
  14 => std_logic_vector'(x"8002618f"),
  15 => std_logic_vector'(x"6050a000"),
  16 => std_logic_vector'(x"63036d00"),
  17 => std_logic_vector'(x"401d0015"),
  18 => std_logic_vector'(x"90002023"),
  19 => std_logic_vector'(x"6d8c6050"),
  20 => std_logic_vector'(x"401e8001"),
  21 => std_logic_vector'(x"90002028"),
  22 => std_logic_vector'(x"618f6043"),
  23 => std_logic_vector'(x"4028800d"),
  24 => std_logic_vector'(x"0028800a"),
  25 => std_logic_vector'(x"00288020"),
  26 => std_logic_vector'(x"608c8020"),
  27 => std_logic_vector'(x"80106011"),
  28 => std_logic_vector'(x"403a6903"),
  29 => std_logic_vector'(x"80086011"),
  30 => std_logic_vector'(x"403e6903"),
  31 => std_logic_vector'(x"80046011"),
  32 => std_logic_vector'(x"40426903"),
  33 => std_logic_vector'(x"6303800f"),
  34 => std_logic_vector'(x"800a6011"),
  35 => std_logic_vector'(x"204a6803"),
  36 => std_logic_vector'(x"004b8030"),
  37 => std_logic_vector'(x"62038037"),
  38 => std_logic_vector'(x"40360028"),
  39 => std_logic_vector'(x"80000032"),
  40 => std_logic_vector'(x"8000608c"),
  41 => std_logic_vector'(x"6127668c"),
  42 => std_logic_vector'(x"6b1d6110"),
  43 => std_logic_vector'(x"6110619c"),
  44 => std_logic_vector'(x"61106127"),
  45 => std_logic_vector'(x"608c6b1d"),
  46 => std_logic_vector'(x"619d6110"),
  47 => std_logic_vector'(x"618f6103"),
  48 => std_logic_vector'(x"20636011"),
  49 => std_logic_vector'(x"608c609d"),
  50 => std_logic_vector'(x"619d6111"),
  51 => std_logic_vector'(x"6000405c"),
  52 => std_logic_vector'(x"62036c00"),
  53 => std_logic_vector'(x"60336110"),
  54 => std_logic_vector'(x"4053618f"),
  55 => std_logic_vector'(x"40536127"),
  56 => std_logic_vector'(x"608c6b1d"),
  57 => std_logic_vector'(x"61276127"),
  58 => std_logic_vector'(x"6b1d4064"),
  59 => std_logic_vector'(x"006d6b1d"),
  60 => std_logic_vector'(x"207c6811"),
  61 => std_logic_vector'(x"007d6103"),
  62 => std_logic_vector'(x"608c608f"),
  63 => std_logic_vector'(x"20826811"),
  64 => std_logic_vector'(x"00836003"),
  65 => std_logic_vector'(x"608c618f"),
  66 => std_logic_vector'(x"61106c11"),
  67 => std_logic_vector'(x"6a038003"),
  68 => std_logic_vector'(x"80ff6903"),
  69 => std_logic_vector'(x"8010638f"),
  70 => std_logic_vector'(x"80106903"),
  71 => std_logic_vector'(x"80106a8f"),
  72 => std_logic_vector'(x"80106a03"),
  73 => std_logic_vector'(x"6c11698f"),
  74 => std_logic_vector'(x"80026110"),
  75 => std_logic_vector'(x"80036303"),
  76 => std_logic_vector'(x"69036a03"),
  77 => std_logic_vector'(x"4093008f"),
  78 => std_logic_vector'(x"800f8001"),
  79 => std_logic_vector'(x"80006a03"),
  80 => std_logic_vector'(x"63006403"),
  81 => std_logic_vector'(x"800120aa"),
  82 => std_logic_vector'(x"6a03800f"),
  83 => std_logic_vector'(x"6403ffff"),
  84 => std_logic_vector'(x"628f6600"),
  85 => std_logic_vector'(x"6024608c"),
  86 => std_logic_vector'(x"63038002"),
  87 => std_logic_vector'(x"801020b6"),
  88 => std_logic_vector'(x"6b116a03"),
  89 => std_logic_vector'(x"6c006000"),
  90 => std_logic_vector'(x"00bb408f"),
  91 => std_logic_vector'(x"6b11408f"),
  92 => std_logic_vector'(x"6c006000"),
  93 => std_logic_vector'(x"6403408b"),
  94 => std_logic_vector'(x"60336b1d"),
  95 => std_logic_vector'(x"405c618f"),
  96 => std_logic_vector'(x"62034093"),
  97 => std_logic_vector'(x"00ab6110"),
  98 => std_logic_vector'(x"80016024"),
  99 => std_logic_vector'(x"20cc6303"),
  100 => std_logic_vector'(x"6a038008"),
  101 => std_logic_vector'(x"00d380ff"),
  102 => std_logic_vector'(x"630380ff"),
  103 => std_logic_vector'(x"800f8001"),
  104 => std_logic_vector'(x"ff006a03"),
  105 => std_logic_vector'(x"6b116403"),
  106 => std_logic_vector'(x"63034093"),
  107 => std_logic_vector'(x"6b1d6403"),
  108 => std_logic_vector'(x"601100ab"),
  109 => std_logic_vector'(x"61104002"),
  110 => std_logic_vector'(x"61110084"),
  111 => std_logic_vector'(x"619c6203"),
  112 => std_logic_vector'(x"651140dd"),
  113 => std_logic_vector'(x"601120e8"),
  114 => std_logic_vector'(x"40284084"),
  115 => std_logic_vector'(x"00e14002"),
  116 => std_logic_vector'(x"c16c005e"),
  117 => std_logic_vector'(x"c168608c"),
  118 => std_logic_vector'(x"c18c608c"),
  119 => std_logic_vector'(x"c160608c"),
  120 => std_logic_vector'(x"c188608c"),
  121 => std_logic_vector'(x"c164608c"),
  122 => std_logic_vector'(x"c19c608c"),
  123 => std_logic_vector'(x"4093608c"),
  124 => std_logic_vector'(x"66008001"),
  125 => std_logic_vector'(x"c164638f"),
  126 => std_logic_vector'(x"60114093"),
  127 => std_logic_vector'(x"60112107"),
  128 => std_logic_vector'(x"62038002"),
  129 => std_logic_vector'(x"40e040d9"),
  130 => std_logic_vector'(x"40f74032"),
  131 => std_logic_vector'(x"618f00fd"),
  132 => std_logic_vector'(x"00026600"),
  133 => std_logic_vector'(x"628f4108"),
  134 => std_logic_vector'(x"40116011"),
  135 => std_logic_vector'(x"01082110"),
  136 => std_logic_vector'(x"8001608c"),
  137 => std_logic_vector'(x"60116a8f"),
  138 => std_logic_vector'(x"211b4011"),
  139 => std_logic_vector'(x"80016600"),
  140 => std_logic_vector'(x"66006903"),
  141 => std_logic_vector'(x"8001011d"),
  142 => std_logic_vector'(x"608c698f"),
  143 => std_logic_vector'(x"6000c16c"),
  144 => std_logic_vector'(x"6e116c8c"),
  145 => std_logic_vector'(x"638f801f"),
  146 => std_logic_vector'(x"61276011"),
  147 => std_logic_vector'(x"6110410a"),
  148 => std_logic_vector'(x"62036b1d"),
  149 => std_logic_vector'(x"8003619c"),
  150 => std_logic_vector'(x"80036203"),
  151 => std_logic_vector'(x"638f6600"),
  152 => std_logic_vector'(x"62034053"),
  153 => std_logic_vector'(x"62006127"),
  154 => std_logic_vector'(x"61116110"),
  155 => std_logic_vector'(x"6f036110"),
  156 => std_logic_vector'(x"6b1d213c"),
  157 => std_logic_vector'(x"013d4002"),
  158 => std_logic_vector'(x"608c6b1d"),
  159 => std_logic_vector'(x"61106600"),
  160 => std_logic_vector'(x"61106600"),
  161 => std_logic_vector'(x"80008001"),
  162 => std_logic_vector'(x"60110130"),
  163 => std_logic_vector'(x"21494011"),
  164 => std_logic_vector'(x"608c013e"),
  165 => std_logic_vector'(x"00116011"),
  166 => std_logic_vector'(x"40096011"),
  167 => std_logic_vector'(x"6c006000"),
  168 => std_logic_vector'(x"60006110"),
  169 => std_logic_vector'(x"405c6c8c"),
  170 => std_logic_vector'(x"61036033"),
  171 => std_logic_vector'(x"60334009"),
  172 => std_logic_vector'(x"6127618f"),
  173 => std_logic_vector'(x"406d6127"),
  174 => std_logic_vector'(x"6b1d6b1d"),
  175 => std_logic_vector'(x"618f006d"),
  176 => std_logic_vector'(x"40536127"),
  177 => std_logic_vector'(x"61106703"),
  178 => std_logic_vector'(x"67036b1d"),
  179 => std_logic_vector'(x"4053638f"),
  180 => std_logic_vector'(x"67034064"),
  181 => std_logic_vector'(x"405e216e"),
  182 => std_logic_vector'(x"01716f03"),
  183 => std_logic_vector'(x"6003400f"),
  184 => std_logic_vector'(x"608c608f"),
  185 => std_logic_vector'(x"40644053"),
  186 => std_logic_vector'(x"21796703"),
  187 => std_logic_vector'(x"6f03405e"),
  188 => std_logic_vector'(x"4017017c"),
  189 => std_logic_vector'(x"608f6003"),
  190 => std_logic_vector'(x"413e608c"),
  191 => std_logic_vector'(x"60030130"),
  192 => std_logic_vector'(x"64030011"),
  193 => std_logic_vector'(x"40640007"),
  194 => std_logic_vector'(x"61270130"),
  195 => std_logic_vector'(x"69038001"),
  196 => std_logic_vector'(x"801f6b11"),
  197 => std_logic_vector'(x"64036a03"),
  198 => std_logic_vector'(x"01136b1d"),
  199 => std_logic_vector'(x"4190418f"),
  200 => std_logic_vector'(x"41924191"),
  201 => std_logic_vector'(x"61274193"),
  202 => std_logic_vector'(x"6a038001"),
  203 => std_logic_vector'(x"801f6111"),
  204 => std_logic_vector'(x"62036903"),
  205 => std_logic_vector'(x"80016110"),
  206 => std_logic_vector'(x"61106a03"),
  207 => std_logic_vector'(x"80006b11"),
  208 => std_logic_vector'(x"21a76803"),
  209 => std_logic_vector'(x"6000c348"),
  210 => std_logic_vector'(x"80006c00"),
  211 => std_logic_vector'(x"6b1d4130"),
  212 => std_logic_vector'(x"6a8f8001"),
  213 => std_logic_vector'(x"6033c348"),
  214 => std_logic_vector'(x"80006103"),
  215 => std_logic_vector'(x"40538000"),
  216 => std_logic_vector'(x"618f418e"),
  217 => std_logic_vector'(x"41b441b3"),
  218 => std_logic_vector'(x"41b641b5"),
  219 => std_logic_vector'(x"612741b7"),
  220 => std_logic_vector'(x"6a038001"),
  221 => std_logic_vector'(x"80006b11"),
  222 => std_logic_vector'(x"21c26803"),
  223 => std_logic_vector'(x"6000c348"),
  224 => std_logic_vector'(x"62036c00"),
  225 => std_logic_vector'(x"80016b1d"),
  226 => std_logic_vector'(x"c3486a8f"),
  227 => std_logic_vector'(x"61036033"),
  228 => std_logic_vector'(x"61108000"),
  229 => std_logic_vector'(x"618f41b2"),
  230 => std_logic_vector'(x"41ce41cd"),
  231 => std_logic_vector'(x"41d041cf"),
  232 => std_logic_vector'(x"612741d1"),
  233 => std_logic_vector'(x"40116011"),
  234 => std_logic_vector'(x"40646127"),
  235 => std_logic_vector'(x"60114130"),
  236 => std_logic_vector'(x"64036b1d"),
  237 => std_logic_vector'(x"6f036b11"),
  238 => std_logic_vector'(x"21e36600"),
  239 => std_logic_vector'(x"410a6b11"),
  240 => std_logic_vector'(x"40026110"),
  241 => std_logic_vector'(x"6b1d6110"),
  242 => std_logic_vector'(x"41cc608c"),
  243 => std_logic_vector'(x"619c6103"),
  244 => std_logic_vector'(x"21f06011"),
  245 => std_logic_vector'(x"40288008"),
  246 => std_logic_vector'(x"40288020"),
  247 => std_logic_vector'(x"40288008"),
  248 => std_logic_vector'(x"40076011"),
  249 => std_logic_vector'(x"608c21f4"),
  250 => std_logic_vector'(x"40644004"),
  251 => std_logic_vector'(x"40846203"),
  252 => std_logic_vector'(x"630380c0"),
  253 => std_logic_vector'(x"400d8080"),
  254 => std_logic_vector'(x"608c21f0"),
  255 => std_logic_vector'(x"6000c19c"),
  256 => std_logic_vector'(x"22046c00"),
  257 => std_logic_vector'(x"4028801e"),
  258 => std_logic_vector'(x"80006127"),
  259 => std_logic_vector'(x"80094023"),
  260 => std_logic_vector'(x"220c6700"),
  261 => std_logic_vector'(x"80206103"),
  262 => std_logic_vector'(x"6700807f"),
  263 => std_logic_vector'(x"61032211"),
  264 => std_logic_vector'(x"60118008"),
  265 => std_logic_vector'(x"4017801f"),
  266 => std_logic_vector'(x"61112228"),
  267 => std_logic_vector'(x"6f036b11"),
  268 => std_logic_vector'(x"c19c2228"),
  269 => std_logic_vector'(x"6c006000"),
  270 => std_logic_vector'(x"22204007"),
  271 => std_logic_vector'(x"40286011"),
  272 => std_logic_vector'(x"40646127"),
  273 => std_logic_vector'(x"6b116203"),
  274 => std_logic_vector'(x"40c46110"),
  275 => std_logic_vector'(x"6b1d4002"),
  276 => std_logic_vector'(x"67008008"),
  277 => std_logic_vector'(x"6127222e"),
  278 => std_logic_vector'(x"6b1d41e8"),
  279 => std_logic_vector'(x"6700800a"),
  280 => std_logic_vector'(x"800d6110"),
  281 => std_logic_vector'(x"64036703"),
  282 => std_logic_vector'(x"600c2206"),
  283 => std_logic_vector'(x"00326003"),
  284 => std_logic_vector'(x"61116127"),
  285 => std_logic_vector'(x"619c6b1d"),
  286 => std_logic_vector'(x"42384238"),
  287 => std_logic_vector'(x"80400238"),
  288 => std_logic_vector'(x"68036111"),
  289 => std_logic_vector'(x"805b6111"),
  290 => std_logic_vector'(x"63036803"),
  291 => std_logic_vector'(x"63038020"),
  292 => std_logic_vector'(x"6511628f"),
  293 => std_logic_vector'(x"6303801f"),
  294 => std_logic_vector'(x"6103224f"),
  295 => std_logic_vector'(x"423f608c"),
  296 => std_logic_vector'(x"423f6110"),
  297 => std_logic_vector'(x"4064658f"),
  298 => std_logic_vector'(x"62038002"),
  299 => std_logic_vector'(x"67034084"),
  300 => std_logic_vector'(x"423c2273"),
  301 => std_logic_vector'(x"62038003"),
  302 => std_logic_vector'(x"40dd6127"),
  303 => std_logic_vector'(x"226f6511"),
  304 => std_logic_vector'(x"40846011"),
  305 => std_logic_vector'(x"40846b11"),
  306 => std_logic_vector'(x"226a4249"),
  307 => std_logic_vector'(x"600c405e"),
  308 => std_logic_vector'(x"608c404f"),
  309 => std_logic_vector'(x"6b1d4002"),
  310 => std_logic_vector'(x"61274002"),
  311 => std_logic_vector'(x"405e025e"),
  312 => std_logic_vector'(x"4051600c"),
  313 => std_logic_vector'(x"004f0274"),
  314 => std_logic_vector'(x"4002608c"),
  315 => std_logic_vector'(x"66008001"),
  316 => std_logic_vector'(x"8002638f"),
  317 => std_logic_vector'(x"40d96203"),
  318 => std_logic_vector'(x"42756203"),
  319 => std_logic_vector'(x"c16c0093"),
  320 => std_logic_vector'(x"6c006000"),
  321 => std_logic_vector'(x"c16c4275"),
  322 => std_logic_vector'(x"618f6033"),
  323 => std_logic_vector'(x"80014093"),
  324 => std_logic_vector'(x"41116303"),
  325 => std_logic_vector'(x"c1640004"),
  326 => std_logic_vector'(x"60114093"),
  327 => std_logic_vector'(x"4253229a"),
  328 => std_logic_vector'(x"60032298"),
  329 => std_logic_vector'(x"60116003"),
  330 => std_logic_vector'(x"61104279"),
  331 => std_logic_vector'(x"608c4286"),
  332 => std_logic_vector'(x"028d40f7"),
  333 => std_logic_vector'(x"423f608c"),
  334 => std_logic_vector'(x"80396011"),
  335 => std_logic_vector'(x"8100400f"),
  336 => std_logic_vector'(x"62036303"),
  337 => std_logic_vector'(x"81606011"),
  338 => std_logic_vector'(x"8127400f"),
  339 => std_logic_vector'(x"410a6303"),
  340 => std_logic_vector'(x"410a8030"),
  341 => std_logic_vector'(x"c1606011"),
  342 => std_logic_vector'(x"6c006000"),
  343 => std_logic_vector'(x"405c6f8f"),
  344 => std_logic_vector'(x"612741c5"),
  345 => std_logic_vector'(x"6b1d41aa"),
  346 => std_logic_vector'(x"6011628f"),
  347 => std_logic_vector'(x"611122cb"),
  348 => std_logic_vector'(x"429b4084"),
  349 => std_logic_vector'(x"22be4007"),
  350 => std_logic_vector'(x"608c6103"),
  351 => std_logic_vector'(x"406d6127"),
  352 => std_logic_vector'(x"6000c160"),
  353 => std_logic_vector'(x"42af6c00"),
  354 => std_logic_vector'(x"414a6b1d"),
  355 => std_logic_vector'(x"406d4130"),
  356 => std_logic_vector'(x"41248001"),
  357 => std_logic_vector'(x"608c02b5"),
  358 => std_logic_vector'(x"40dd6127"),
  359 => std_logic_vector'(x"22d56511"),
  360 => std_logic_vector'(x"61116b11"),
  361 => std_logic_vector'(x"400240c4"),
  362 => std_logic_vector'(x"6b1d02ce"),
  363 => std_logic_vector'(x"005e6103"),
  364 => std_logic_vector'(x"405340dd"),
  365 => std_logic_vector'(x"65116127"),
  366 => std_logic_vector'(x"6b1122e6"),
  367 => std_logic_vector'(x"61114084"),
  368 => std_logic_vector'(x"6b1d40c4"),
  369 => std_logic_vector'(x"61274002"),
  370 => std_logic_vector'(x"02db4002"),
  371 => std_logic_vector'(x"005e600c"),
  372 => std_logic_vector'(x"22f66011"),
  373 => std_logic_vector'(x"61274004"),
  374 => std_logic_vector'(x"6b116111"),
  375 => std_logic_vector'(x"40846203"),
  376 => std_logic_vector'(x"6b116111"),
  377 => std_logic_vector'(x"40c46203"),
  378 => std_logic_vector'(x"02e86b1d"),
  379 => std_logic_vector'(x"005e6103"),
  380 => std_logic_vector'(x"608c6127"),
  381 => std_logic_vector'(x"014cc17c"),
  382 => std_logic_vector'(x"0153c17c"),
  383 => std_logic_vector'(x"6000c184"),
  384 => std_logic_vector'(x"80216c8c"),
  385 => std_logic_vector'(x"43016f8f"),
  386 => std_logic_vector'(x"61270007"),
  387 => std_logic_vector'(x"40846111"),
  388 => std_logic_vector'(x"42f86b11"),
  389 => std_logic_vector'(x"230f6300"),
  390 => std_logic_vector'(x"41248001"),
  391 => std_logic_vector'(x"6b1d0306"),
  392 => std_logic_vector'(x"42fa618f"),
  393 => std_logic_vector'(x"6000c188"),
  394 => std_logic_vector'(x"41246c00"),
  395 => std_logic_vector'(x"43058602"),
  396 => std_logic_vector'(x"61276111"),
  397 => std_logic_vector'(x"43058606"),
  398 => std_logic_vector'(x"80014064"),
  399 => std_logic_vector'(x"62034078"),
  400 => std_logic_vector'(x"610342fa"),
  401 => std_logic_vector'(x"c188410a"),
  402 => std_logic_vector'(x"61036033"),
  403 => std_logic_vector'(x"6b1d6103"),
  404 => std_logic_vector'(x"010a405c"),
  405 => std_logic_vector'(x"6000c190"),
  406 => std_logic_vector'(x"000d6c00"),
  407 => std_logic_vector'(x"6033c190"),
  408 => std_logic_vector'(x"42fa6103"),
  409 => std_logic_vector'(x"6000c188"),
  410 => std_logic_vector'(x"41246c00"),
  411 => std_logic_vector'(x"61276111"),
  412 => std_logic_vector'(x"43058654"),
  413 => std_logic_vector'(x"80014064"),
  414 => std_logic_vector'(x"62034078"),
  415 => std_logic_vector'(x"610342fa"),
  416 => std_logic_vector'(x"c188410a"),
  417 => std_logic_vector'(x"61036033"),
  418 => std_logic_vector'(x"6b1d6103"),
  419 => std_logic_vector'(x"010a405c"),
  420 => std_logic_vector'(x"0066c16c"),
  421 => std_logic_vector'(x"6033411e"),
  422 => std_logic_vector'(x"80046103"),
  423 => std_logic_vector'(x"411e0348"),
  424 => std_logic_vector'(x"800240ab"),
  425 => std_logic_vector'(x"411e0348"),
  426 => std_logic_vector'(x"800140c4"),
  427 => std_logic_vector'(x"c1680348"),
  428 => std_logic_vector'(x"6c006000"),
  429 => std_logic_vector'(x"800240ab"),
  430 => std_logic_vector'(x"0066c168"),
  431 => std_logic_vector'(x"6000c170"),
  432 => std_logic_vector'(x"40606c00"),
  433 => std_logic_vector'(x"c1642366"),
  434 => std_logic_vector'(x"618f6033"),
  435 => std_logic_vector'(x"c168608c"),
  436 => std_logic_vector'(x"6c006000"),
  437 => std_logic_vector'(x"6033c178"),
  438 => std_logic_vector'(x"6011618f"),
  439 => std_logic_vector'(x"40dd4353"),
  440 => std_logic_vector'(x"23756511"),
  441 => std_logic_vector'(x"435340d9"),
  442 => std_logic_vector'(x"005e0370"),
  443 => std_logic_vector'(x"411e427f"),
  444 => std_logic_vector'(x"6033c170"),
  445 => std_logic_vector'(x"c1646103"),
  446 => std_logic_vector'(x"6c006000"),
  447 => std_logic_vector'(x"4311434f"),
  448 => std_logic_vector'(x"427f436d"),
  449 => std_logic_vector'(x"6000c168"),
  450 => std_logic_vector'(x"434f6c00"),
  451 => std_logic_vector'(x"6000c168"),
  452 => std_logic_vector'(x"c1746c00"),
  453 => std_logic_vector'(x"61036033"),
  454 => std_logic_vector'(x"c1700367"),
  455 => std_logic_vector'(x"6c006000"),
  456 => std_logic_vector'(x"40936011"),
  457 => std_logic_vector'(x"64038001"),
  458 => std_logic_vector'(x"00ab6110"),
  459 => std_logic_vector'(x"c18c8003"),
  460 => std_logic_vector'(x"618f6033"),
  461 => std_logic_vector'(x"c18c8000"),
  462 => std_logic_vector'(x"618f6033"),
  463 => std_logic_vector'(x"03964376"),
  464 => std_logic_vector'(x"c168427f"),
  465 => std_logic_vector'(x"6c006000"),
  466 => std_logic_vector'(x"c1746011"),
  467 => std_logic_vector'(x"61036033"),
  468 => std_logic_vector'(x"c1708000"),
  469 => std_logic_vector'(x"61036033"),
  470 => std_logic_vector'(x"03964367"),
  471 => std_logic_vector'(x"60116b1d"),
  472 => std_logic_vector'(x"43574093"),
  473 => std_logic_vector'(x"62038002"),
  474 => std_logic_vector'(x"608c6127"),
  475 => std_logic_vector'(x"6000c168"),
  476 => std_logic_vector'(x"80016c00"),
  477 => std_logic_vector'(x"628f6600"),
  478 => std_logic_vector'(x"6b1d6103"),
  479 => std_logic_vector'(x"c1946b1d"),
  480 => std_logic_vector'(x"61036033"),
  481 => std_logic_vector'(x"608c6127"),
  482 => std_logic_vector'(x"80016011"),
  483 => std_logic_vector'(x"6a03800f"),
  484 => std_logic_vector'(x"6403e000"),
  485 => std_logic_vector'(x"c0006303"),
  486 => std_logic_vector'(x"61106703"),
  487 => std_logic_vector'(x"63039fff"),
  488 => std_logic_vector'(x"87784111"),
  489 => std_logic_vector'(x"638f400d"),
  490 => std_logic_vector'(x"6000c168"),
  491 => std_logic_vector'(x"c1746c00"),
  492 => std_logic_vector'(x"6c006000"),
  493 => std_logic_vector'(x"23e9400d"),
  494 => std_logic_vector'(x"409343b6"),
  495 => std_logic_vector'(x"23e943c4"),
  496 => std_logic_vector'(x"409343b6"),
  497 => std_logic_vector'(x"6503c000"),
  498 => std_logic_vector'(x"40ab43b6"),
  499 => std_logic_vector'(x"608c43ae"),
  500 => std_logic_vector'(x"43ae608c"),
  501 => std_logic_vector'(x"608c608c"),
  502 => std_logic_vector'(x"43d4435e"),
  503 => std_logic_vector'(x"c168039a"),
  504 => std_logic_vector'(x"6c006000"),
  505 => std_logic_vector'(x"0357a000"),
  506 => std_logic_vector'(x"6000c168"),
  507 => std_logic_vector'(x"80006c00"),
  508 => std_logic_vector'(x"60110357"),
  509 => std_logic_vector'(x"c1684093"),
  510 => std_logic_vector'(x"6c006000"),
  511 => std_logic_vector'(x"64034113"),
  512 => std_logic_vector'(x"40ab6110"),
  513 => std_logic_vector'(x"c1680367"),
  514 => std_logic_vector'(x"6c006000"),
  515 => std_logic_vector'(x"03570113"),
  516 => std_logic_vector'(x"6403a000"),
  517 => std_logic_vector'(x"80010357"),
  518 => std_logic_vector'(x"6a03800f"),
  519 => std_logic_vector'(x"6403e080"),
  520 => std_logic_vector'(x"e0806303"),
  521 => std_logic_vector'(x"6011678f"),
  522 => std_logic_vector'(x"80014093"),
  523 => std_logic_vector'(x"6a03800f"),
  524 => std_logic_vector'(x"64038000"),
  525 => std_logic_vector'(x"40156303"),
  526 => std_logic_vector'(x"80026110"),
  527 => std_logic_vector'(x"40936203"),
  528 => std_logic_vector'(x"6703e08c"),
  529 => std_logic_vector'(x"6011638f"),
  530 => std_logic_vector'(x"440b4093"),
  531 => std_logic_vector'(x"40932430"),
  532 => std_logic_vector'(x"800f8001"),
  533 => std_logic_vector'(x"ff736a03"),
  534 => std_logic_vector'(x"63036403"),
  535 => std_logic_vector'(x"043a4357"),
  536 => std_logic_vector'(x"44136011"),
  537 => std_logic_vector'(x"40932436"),
  538 => std_logic_vector'(x"043a4357"),
  539 => std_logic_vector'(x"c0004113"),
  540 => std_logic_vector'(x"03576403"),
  541 => std_logic_vector'(x"6b1d608c"),
  542 => std_logic_vector'(x"c1704113"),
  543 => std_logic_vector'(x"6c006000"),
  544 => std_logic_vector'(x"80024279"),
  545 => std_logic_vector'(x"00ab6203"),
  546 => std_logic_vector'(x"6000c174"),
  547 => std_logic_vector'(x"04236c00"),
  548 => std_logic_vector'(x"c1946b1d"),
  549 => std_logic_vector'(x"6c006000"),
  550 => std_logic_vector'(x"61276127"),
  551 => std_logic_vector'(x"c1946111"),
  552 => std_logic_vector'(x"61036033"),
  553 => std_logic_vector'(x"010a6110"),
  554 => std_logic_vector'(x"c1946b1d"),
  555 => std_logic_vector'(x"6c006000"),
  556 => std_logic_vector'(x"61276127"),
  557 => std_logic_vector'(x"c1946111"),
  558 => std_logic_vector'(x"61036033"),
  559 => std_logic_vector'(x"410a6110"),
  560 => std_logic_vector'(x"00076011"),
  561 => std_logic_vector'(x"62038001"),
  562 => std_logic_vector'(x"c198609d"),
  563 => std_logic_vector'(x"6c006000"),
  564 => std_logic_vector'(x"c1988000"),
  565 => std_logic_vector'(x"61036033"),
  566 => std_logic_vector'(x"44238890"),
  567 => std_logic_vector'(x"43ae4403"),
  568 => std_logic_vector'(x"608c6127"),
  569 => std_logic_vector'(x"6000c198"),
  570 => std_logic_vector'(x"60116c00"),
  571 => std_logic_vector'(x"60112481"),
  572 => std_logic_vector'(x"61104093"),
  573 => std_logic_vector'(x"6000c168"),
  574 => std_logic_vector'(x"41136c00"),
  575 => std_logic_vector'(x"40ab6110"),
  576 => std_logic_vector'(x"61030475"),
  577 => std_logic_vector'(x"6033c198"),
  578 => std_logic_vector'(x"87786103"),
  579 => std_logic_vector'(x"43ae0423"),
  580 => std_logic_vector'(x"88c46b1d"),
  581 => std_logic_vector'(x"43ef4423"),
  582 => std_logic_vector'(x"44076110"),
  583 => std_logic_vector'(x"047243f9"),
  584 => std_logic_vector'(x"40116111"),
  585 => std_logic_vector'(x"60242499"),
  586 => std_logic_vector'(x"6b1d6203"),
  587 => std_logic_vector'(x"6f036111"),
  588 => std_logic_vector'(x"6024049e"),
  589 => std_logic_vector'(x"6b1d6203"),
  590 => std_logic_vector'(x"00176111"),
  591 => std_logic_vector'(x"43ae608c"),
  592 => std_logic_vector'(x"89206b1d"),
  593 => std_logic_vector'(x"44084423"),
  594 => std_logic_vector'(x"43ae0472"),
  595 => std_logic_vector'(x"c1686b1d"),
  596 => std_logic_vector'(x"6c006000"),
  597 => std_logic_vector'(x"6000c198"),
  598 => std_logic_vector'(x"43576c00"),
  599 => std_logic_vector'(x"6033c198"),
  600 => std_logic_vector'(x"c198618f"),
  601 => std_logic_vector'(x"6c006000"),
  602 => std_logic_vector'(x"c1988000"),
  603 => std_logic_vector'(x"61036033"),
  604 => std_logic_vector'(x"442388a8"),
  605 => std_logic_vector'(x"c16843ef"),
  606 => std_logic_vector'(x"6c006000"),
  607 => std_logic_vector'(x"6000c198"),
  608 => std_logic_vector'(x"43576c00"),
  609 => std_logic_vector'(x"6033c198"),
  610 => std_logic_vector'(x"43f96103"),
  611 => std_logic_vector'(x"43ae4403"),
  612 => std_logic_vector'(x"608c6127"),
  613 => std_logic_vector'(x"6b116b1d"),
  614 => std_logic_vector'(x"6000c194"),
  615 => std_logic_vector'(x"62036c00"),
  616 => std_logic_vector'(x"61276110"),
  617 => std_logic_vector'(x"6b1d608c"),
  618 => std_logic_vector'(x"6b1d6b1d"),
  619 => std_logic_vector'(x"40646b1d"),
  620 => std_logic_vector'(x"40576203"),
  621 => std_logic_vector'(x"61276127"),
  622 => std_logic_vector'(x"61274057"),
  623 => std_logic_vector'(x"608c6127"),
  624 => std_logic_vector'(x"6b1d43ae"),
  625 => std_logic_vector'(x"04238778"),
  626 => std_logic_vector'(x"c160800a"),
  627 => std_logic_vector'(x"618f6033"),
  628 => std_logic_vector'(x"618f6033"),
  629 => std_logic_vector'(x"658f628f"),
  630 => std_logic_vector'(x"648f638f"),
  631 => std_logic_vector'(x"678f668c"),
  632 => std_logic_vector'(x"6f8f688f"),
  633 => std_logic_vector'(x"609d619c"),
  634 => std_logic_vector'(x"619d618f"),
  635 => std_logic_vector'(x"6000608f"),
  636 => std_logic_vector'(x"60436c8c"),
  637 => std_logic_vector'(x"6050618f"),
  638 => std_logic_vector'(x"698f6d8c"),
  639 => std_logic_vector'(x"43ae6a8f"),
  640 => std_logic_vector'(x"608c6127"),
  641 => std_logic_vector'(x"6b1d43ae"),
  642 => std_logic_vector'(x"43ae608c"),
  643 => std_logic_vector'(x"608c6b11"),
  644 => std_logic_vector'(x"62036b1d"),
  645 => std_logic_vector'(x"608c6127"),
  646 => std_logic_vector'(x"251e4060"),
  647 => std_logic_vector'(x"40288065"),
  648 => std_logic_vector'(x"40288072"),
  649 => std_logic_vector'(x"40288072"),
  650 => std_logic_vector'(x"4028806f"),
  651 => std_logic_vector'(x"40288072"),
  652 => std_logic_vector'(x"4028803a"),
  653 => std_logic_vector'(x"404d4032"),
  654 => std_logic_vector'(x"02f88002"),
  655 => std_logic_vector'(x"4108608c"),
  656 => std_logic_vector'(x"050c6303"),
  657 => std_logic_vector'(x"45246110"),
  658 => std_logic_vector'(x"40116011"),
  659 => std_logic_vector'(x"6600252c"),
  660 => std_logic_vector'(x"43ae4524"),
  661 => std_logic_vector'(x"05466600"),
  662 => std_logic_vector'(x"ffff6011"),
  663 => std_logic_vector'(x"63036600"),
  664 => std_logic_vector'(x"6011253f"),
  665 => std_logic_vector'(x"6903800f"),
  666 => std_logic_vector'(x"800f4524"),
  667 => std_logic_vector'(x"43ae4524"),
  668 => std_logic_vector'(x"ffff6a03"),
  669 => std_logic_vector'(x"45246303"),
  670 => std_logic_vector'(x"640343ae"),
  671 => std_logic_vector'(x"80010546"),
  672 => std_logic_vector'(x"6a03800f"),
  673 => std_logic_vector'(x"64038000"),
  674 => std_logic_vector'(x"03576403"),
  675 => std_logic_vector'(x"6003608c"),
  676 => std_logic_vector'(x"800d4015"),
  677 => std_logic_vector'(x"6127051f"),
  678 => std_logic_vector'(x"40846111"),
  679 => std_logic_vector'(x"67036b1d"),
  680 => std_logic_vector'(x"40156111"),
  681 => std_logic_vector'(x"60246303"),
  682 => std_logic_vector'(x"63038001"),
  683 => std_logic_vector'(x"6b1d4124"),
  684 => std_logic_vector'(x"8000608c"),
  685 => std_logic_vector'(x"406d8000"),
  686 => std_logic_vector'(x"454b802d"),
  687 => std_logic_vector'(x"42b56127"),
  688 => std_logic_vector'(x"454b802e"),
  689 => std_logic_vector'(x"45472569"),
  690 => std_logic_vector'(x"25676b1d"),
  691 => std_logic_vector'(x"8a44413e"),
  692 => std_logic_vector'(x"4547608c"),
  693 => std_logic_vector'(x"6b1d6103"),
  694 => std_logic_vector'(x"4108256e"),
  695 => std_logic_vector'(x"608c8a48"),
  696 => std_logic_vector'(x"6000c160"),
  697 => std_logic_vector'(x"61276c00"),
  698 => std_logic_vector'(x"455944e5"),
  699 => std_logic_vector'(x"04e56b1d"),
  700 => std_logic_vector'(x"67038003"),
  701 => std_logic_vector'(x"40846111"),
  702 => std_logic_vector'(x"67038027"),
  703 => std_logic_vector'(x"61106303"),
  704 => std_logic_vector'(x"40024002"),
  705 => std_logic_vector'(x"80274084"),
  706 => std_logic_vector'(x"638f6703"),
  707 => std_logic_vector'(x"454b8024"),
  708 => std_logic_vector'(x"8010258c"),
  709 => std_logic_vector'(x"608c4570"),
  710 => std_logic_vector'(x"454b8023"),
  711 => std_logic_vector'(x"800a2592"),
  712 => std_logic_vector'(x"608c4570"),
  713 => std_logic_vector'(x"454b8025"),
  714 => std_logic_vector'(x"80022598"),
  715 => std_logic_vector'(x"608c4570"),
  716 => std_logic_vector'(x"45784064"),
  717 => std_logic_vector'(x"610325a0"),
  718 => std_logic_vector'(x"40844002"),
  719 => std_logic_vector'(x"608c456e"),
  720 => std_logic_vector'(x"45860559"),
  721 => std_logic_vector'(x"4311618f"),
  722 => std_logic_vector'(x"6011428b"),
  723 => std_logic_vector'(x"800d4007"),
  724 => std_logic_vector'(x"4011451f"),
  725 => std_logic_vector'(x"452425ad"),
  726 => std_logic_vector'(x"04238846"),
  727 => std_logic_vector'(x"02f84586"),
  728 => std_logic_vector'(x"02f84508"),
  729 => std_logic_vector'(x"02f805a1"),
  730 => std_logic_vector'(x"05ae0423"),
  731 => std_logic_vector'(x"431102f8"),
  732 => std_logic_vector'(x"25c36011"),
  733 => std_logic_vector'(x"c18c428b"),
  734 => std_logic_vector'(x"6c006000"),
  735 => std_logic_vector'(x"40026203"),
  736 => std_logic_vector'(x"45b04111"),
  737 => std_logic_vector'(x"005e05b7"),
  738 => std_logic_vector'(x"400742fe"),
  739 => std_logic_vector'(x"25d16011"),
  740 => std_logic_vector'(x"6011c1a0"),
  741 => std_logic_vector'(x"41fe8080"),
  742 => std_logic_vector'(x"800042fc"),
  743 => std_logic_vector'(x"6033c188"),
  744 => std_logic_vector'(x"608c618f"),
  745 => std_logic_vector'(x"612742fa"),
  746 => std_logic_vector'(x"c1886127"),
  747 => std_logic_vector'(x"6c006000"),
  748 => std_logic_vector'(x"42fe6127"),
  749 => std_logic_vector'(x"80006127"),
  750 => std_logic_vector'(x"c1846600"),
  751 => std_logic_vector'(x"61036033"),
  752 => std_logic_vector'(x"800042fc"),
  753 => std_logic_vector'(x"6033c188"),
  754 => std_logic_vector'(x"45b76103"),
  755 => std_logic_vector'(x"c1846b1d"),
  756 => std_logic_vector'(x"61036033"),
  757 => std_logic_vector'(x"c1886b1d"),
  758 => std_logic_vector'(x"61036033"),
  759 => std_logic_vector'(x"6b1d6b1d"),
  760 => std_logic_vector'(x"45c402fc"),
  761 => std_logic_vector'(x"45b76103"),
  762 => std_logic_vector'(x"806f4032"),
  763 => std_logic_vector'(x"806b4028"),
  764 => std_logic_vector'(x"402e4028"),
  765 => std_logic_vector'(x"608c05f1"),
  766 => std_logic_vector'(x"c19c44e4"),
  767 => std_logic_vector'(x"c15c4019"),
  768 => std_logic_vector'(x"428b8004"),
  769 => std_logic_vector'(x"42f82605"),
  770 => std_logic_vector'(x"405e0606"),
  771 => std_logic_vector'(x"42fa05f1"),
  772 => std_logic_vector'(x"c1886003"),
  773 => std_logic_vector'(x"608c04e8"),
  774 => std_logic_vector'(x"608c0002"),
  775 => std_logic_vector'(x"8000608c"),
  776 => std_logic_vector'(x"050c6600"),
  777 => std_logic_vector'(x"4311608c"),
  778 => std_logic_vector'(x"4007428b"),
  779 => std_logic_vector'(x"6600800c"),
  780 => std_logic_vector'(x"050c6303"),
  781 => std_logic_vector'(x"4613608c"),
  782 => std_logic_vector'(x"608c0524"),
  783 => std_logic_vector'(x"61034311"),
  784 => std_logic_vector'(x"608c0084"),
  785 => std_logic_vector'(x"0524461e"),
  786 => std_logic_vector'(x"8029608c"),
  787 => std_logic_vector'(x"005e432e"),
  788 => std_logic_vector'(x"43f4608c"),
  789 => std_logic_vector'(x"03f96110"),
  790 => std_logic_vector'(x"43ef608c"),
  791 => std_logic_vector'(x"608c6110"),
  792 => std_logic_vector'(x"03f94407"),
  793 => std_logic_vector'(x"411e608c"),
  794 => std_logic_vector'(x"c16c412b"),
  795 => std_logic_vector'(x"608c04e8"),
  796 => std_logic_vector'(x"40576b1d"),
  797 => std_logic_vector'(x"61276110"),
  798 => std_logic_vector'(x"61276127"),
  799 => std_logic_vector'(x"4502608c"),
  800 => std_logic_vector'(x"89e44502"),
  801 => std_logic_vector'(x"608c0423"),
  802 => std_logic_vector'(x"6b1d6b1d"),
  803 => std_logic_vector'(x"61106b1d"),
  804 => std_logic_vector'(x"46384064"),
  805 => std_logic_vector'(x"61274053"),
  806 => std_logic_vector'(x"439e608c"),
  807 => std_logic_vector'(x"411e4633"),
  808 => std_logic_vector'(x"03ec4524"),
  809 => std_logic_vector'(x"4093608c"),
  810 => std_logic_vector'(x"6303ffff"),
  811 => std_logic_vector'(x"464d608c"),
  812 => std_logic_vector'(x"400b8002"),
  813 => std_logic_vector'(x"608c0348"),
  814 => std_logic_vector'(x"434a464d"),
  815 => std_logic_vector'(x"443b434a"),
  816 => std_logic_vector'(x"608c014c"),
  817 => std_logic_vector'(x"40724072"),
  818 => std_logic_vector'(x"26674167"),
  819 => std_logic_vector'(x"005e406d"),
  820 => std_logic_vector'(x"4072608c"),
  821 => std_logic_vector'(x"41674072"),
  822 => std_logic_vector'(x"266f6600"),
  823 => std_logic_vector'(x"005e406d"),
  824 => std_logic_vector'(x"414a608c"),
  825 => std_logic_vector'(x"608c0130"),
  826 => std_logic_vector'(x"65034064"),
  827 => std_logic_vector'(x"410c6127"),
  828 => std_logic_vector'(x"410c6110"),
  829 => std_logic_vector'(x"6b1d41aa"),
  830 => std_logic_vector'(x"267f4011"),
  831 => std_logic_vector'(x"608c013e"),
  832 => std_logic_vector'(x"40646127"),
  833 => std_logic_vector'(x"60116403"),
  834 => std_logic_vector'(x"61032688"),
  835 => std_logic_vector'(x"8001413e"),
  836 => std_logic_vector'(x"62036b1d"),
  837 => std_logic_vector'(x"608c0108"),
  838 => std_logic_vector'(x"65034064"),
  839 => std_logic_vector'(x"61276127"),
  840 => std_logic_vector'(x"6b1d4145"),
  841 => std_logic_vector'(x"4638410c"),
  842 => std_logic_vector'(x"41aa6b11"),
  843 => std_logic_vector'(x"6b1d8000"),
  844 => std_logic_vector'(x"61106b1d"),
  845 => std_logic_vector'(x"413041aa"),
  846 => std_logic_vector'(x"40116b1d"),
  847 => std_logic_vector'(x"068026a0"),
  848 => std_logic_vector'(x"6111608c"),
  849 => std_logic_vector'(x"61276127"),
  850 => std_logic_vector'(x"40116011"),
  851 => std_logic_vector'(x"468026a8"),
  852 => std_logic_vector'(x"41e56b11"),
  853 => std_logic_vector'(x"40534053"),
  854 => std_logic_vector'(x"41e56b1d"),
  855 => std_logic_vector'(x"61106003"),
  856 => std_logic_vector'(x"40116b1d"),
  857 => std_logic_vector'(x"013e26b4"),
  858 => std_logic_vector'(x"6127608c"),
  859 => std_logic_vector'(x"6b1d468c"),
  860 => std_logic_vector'(x"608c06a1"),
  861 => std_logic_vector'(x"8000464d"),
  862 => std_logic_vector'(x"608c034a"),
  863 => std_logic_vector'(x"4524439e"),
  864 => std_logic_vector'(x"608c03ec"),
  865 => std_logic_vector'(x"26c54011"),
  866 => std_logic_vector'(x"608c0108"),
  867 => std_logic_vector'(x"65034064"),
  868 => std_logic_vector'(x"61116127"),
  869 => std_logic_vector'(x"410c6127"),
  870 => std_logic_vector'(x"41456127"),
  871 => std_logic_vector'(x"41e56b1d"),
  872 => std_logic_vector'(x"6b1d6110"),
  873 => std_logic_vector'(x"611046c2"),
  874 => std_logic_vector'(x"06c26b1d"),
  875 => std_logic_vector'(x"6011608c"),
  876 => std_logic_vector'(x"40646127"),
  877 => std_logic_vector'(x"61276503"),
  878 => std_logic_vector'(x"41456127"),
  879 => std_logic_vector'(x"410c6b11"),
  880 => std_logic_vector'(x"6b1d41e5"),
  881 => std_logic_vector'(x"26e74011"),
  882 => std_logic_vector'(x"41086110"),
  883 => std_logic_vector'(x"6b1d6110"),
  884 => std_logic_vector'(x"26f24011"),
  885 => std_logic_vector'(x"61114108"),
  886 => std_logic_vector'(x"6b1126f2"),
  887 => std_logic_vector'(x"410a4053"),
  888 => std_logic_vector'(x"40046110"),
  889 => std_logic_vector'(x"61036b1d"),
  890 => std_logic_vector'(x"6127608c"),
  891 => std_logic_vector'(x"6b1d4674"),
  892 => std_logic_vector'(x"608c06c6"),
  893 => std_logic_vector'(x"600346f5"),
  894 => std_logic_vector'(x"6011608c"),
  895 => std_logic_vector'(x"27034013"),
  896 => std_logic_vector'(x"40044032"),
  897 => std_logic_vector'(x"610306fd"),
  898 => std_logic_vector'(x"c798608c"),
  899 => std_logic_vector'(x"c7da608c"),
  900 => std_logic_vector'(x"c7ec608c"),
  901 => std_logic_vector'(x"c7da608c"),
  902 => std_logic_vector'(x"04e8c7ec"),
  903 => std_logic_vector'(x"8000608c"),
  904 => std_logic_vector'(x"c7ec6600"),
  905 => std_logic_vector'(x"c7ec4066"),
  906 => std_logic_vector'(x"00c444f7"),
  907 => std_logic_vector'(x"4011608c"),
  908 => std_logic_vector'(x"802d271b"),
  909 => std_logic_vector'(x"608c070f"),
  910 => std_logic_vector'(x"c1608000"),
  911 => std_logic_vector'(x"41e544f7"),
  912 => std_logic_vector'(x"c1606127"),
  913 => std_logic_vector'(x"41e544f7"),
  914 => std_logic_vector'(x"80096110"),
  915 => std_logic_vector'(x"68036111"),
  916 => std_logic_vector'(x"63038007"),
  917 => std_logic_vector'(x"80306203"),
  918 => std_logic_vector'(x"470f6203"),
  919 => std_logic_vector'(x"608c6b1d"),
  920 => std_logic_vector'(x"4064471c"),
  921 => std_logic_vector'(x"27304181"),
  922 => std_logic_vector'(x"405e608c"),
  923 => std_logic_vector'(x"44f7c7ec"),
  924 => std_logic_vector'(x"6111c7da"),
  925 => std_logic_vector'(x"608c010a"),
  926 => std_logic_vector'(x"60116127"),
  927 => std_logic_vector'(x"41456127"),
  928 => std_logic_vector'(x"4730470b"),
  929 => std_logic_vector'(x"47176b1d"),
  930 => std_logic_vector'(x"6b1d4735"),
  931 => std_logic_vector'(x"410a6111"),
  932 => std_logic_vector'(x"00e046fd"),
  933 => std_logic_vector'(x"8000608c"),
  934 => std_logic_vector'(x"0032473c"),
  935 => std_logic_vector'(x"414a608c"),
  936 => std_logic_vector'(x"608c074b"),
  937 => std_logic_vector'(x"074b8000"),
  938 => std_logic_vector'(x"6127608c"),
  939 => std_logic_vector'(x"6b1d414a"),
  940 => std_logic_vector'(x"608c073c"),
  941 => std_logic_vector'(x"61108000"),
  942 => std_logic_vector'(x"608c073c"),
  943 => std_logic_vector'(x"40646127"),
  944 => std_logic_vector'(x"27656f03"),
  945 => std_logic_vector'(x"42e86b1d"),
  946 => std_logic_vector'(x"6b1d0767"),
  947 => std_logic_vector'(x"608c02d8"),
  948 => std_logic_vector'(x"612742fa"),
  949 => std_logic_vector'(x"44f7c188"),
  950 => std_logic_vector'(x"40846203"),
  951 => std_logic_vector'(x"67036111"),
  952 => std_logic_vector'(x"c1886b1d"),
  953 => std_logic_vector'(x"650344f7"),
  954 => std_logic_vector'(x"277a6303"),
  955 => std_logic_vector'(x"c1888001"),
  956 => std_logic_vector'(x"07684066"),
  957 => std_logic_vector'(x"6011432e"),
  958 => std_logic_vector'(x"40c4c798"),
  959 => std_logic_vector'(x"4002c798"),
  960 => std_logic_vector'(x"42d86110"),
  961 => std_logic_vector'(x"608cc798"),
  962 => std_logic_vector'(x"414a6127"),
  963 => std_logic_vector'(x"06c66b1d"),
  964 => std_logic_vector'(x"4784608c"),
  965 => std_logic_vector'(x"608c6003"),
  966 => std_logic_vector'(x"61034784"),
  967 => std_logic_vector'(x"411e608c"),
  968 => std_logic_vector'(x"80224524"),
  969 => std_logic_vector'(x"036d432e"),
  970 => std_logic_vector'(x"411e608c"),
  971 => std_logic_vector'(x"81b24524"),
  972 => std_logic_vector'(x"036d4423"),
  973 => std_logic_vector'(x"40d9608c"),
  974 => std_logic_vector'(x"608c00e0"),
  975 => std_logic_vector'(x"432e8022"),
  976 => std_logic_vector'(x"44f7c18c"),
  977 => std_logic_vector'(x"411e27a9"),
  978 => std_logic_vector'(x"436d4524"),
  979 => std_logic_vector'(x"44238f36"),
  980 => std_logic_vector'(x"00e007aa"),
  981 => std_logic_vector'(x"c000608c"),
  982 => std_logic_vector'(x"44f7c168"),
  983 => std_logic_vector'(x"8001410a"),
  984 => std_logic_vector'(x"6a03800f"),
  985 => std_logic_vector'(x"64038000"),
  986 => std_logic_vector'(x"410a411e"),
  987 => std_logic_vector'(x"608c6203"),
  988 => std_logic_vector'(x"012b411e"),
  989 => std_logic_vector'(x"4060608c"),
  990 => std_logic_vector'(x"611027c3"),
  991 => std_logic_vector'(x"40046127"),
  992 => std_logic_vector'(x"6b1d47bb"),
  993 => std_logic_vector'(x"608c6110"),
  994 => std_logic_vector'(x"27cd4060"),
  995 => std_logic_vector'(x"61276110"),
  996 => std_logic_vector'(x"47c44004"),
  997 => std_logic_vector'(x"61106b1d"),
  998 => std_logic_vector'(x"601107ce"),
  999 => std_logic_vector'(x"8000608c"),
  1000 => std_logic_vector'(x"608c02cc"),
  1001 => std_logic_vector'(x"410a6111"),
  1002 => std_logic_vector'(x"410a6127"),
  1003 => std_logic_vector'(x"6f036b1d"),
  1004 => std_logic_vector'(x"8029608c"),
  1005 => std_logic_vector'(x"00e0432e"),
  1006 => std_logic_vector'(x"40d9608c"),
  1007 => std_logic_vector'(x"6011428b"),
  1008 => std_logic_vector'(x"27e54007"),
  1009 => std_logic_vector'(x"4004405e"),
  1010 => std_logic_vector'(x"608c8000"),
  1011 => std_logic_vector'(x"04234613"),
  1012 => std_logic_vector'(x"c908608c"),
  1013 => std_logic_vector'(x"8022608c"),
  1014 => std_logic_vector'(x"c18c432e"),
  1015 => std_logic_vector'(x"27f244f7"),
  1016 => std_logic_vector'(x"07f84795"),
  1017 => std_logic_vector'(x"c908405c"),
  1018 => std_logic_vector'(x"42d86110"),
  1019 => std_logic_vector'(x"6110c908"),
  1020 => std_logic_vector'(x"8000608c"),
  1021 => std_logic_vector'(x"4002608c"),
  1022 => std_logic_vector'(x"442389ea"),
  1023 => std_logic_vector'(x"442389de"),
  1024 => std_logic_vector'(x"89e843ef"),
  1025 => std_logic_vector'(x"61104423"),
  1026 => std_logic_vector'(x"6127608c"),
  1027 => std_logic_vector'(x"6b1d4629"),
  1028 => std_logic_vector'(x"89e8608c"),
  1029 => std_logic_vector'(x"60114423"),
  1030 => std_logic_vector'(x"61102811"),
  1031 => std_logic_vector'(x"400443f9"),
  1032 => std_logic_vector'(x"6103080b"),
  1033 => std_logic_vector'(x"8010608c"),
  1034 => std_logic_vector'(x"04e8c160"),
  1035 => std_logic_vector'(x"c188608c"),
  1036 => std_logic_vector'(x"800144f7"),
  1037 => std_logic_vector'(x"6103608c"),
  1038 => std_logic_vector'(x"44e8c188"),
  1039 => std_logic_vector'(x"608c0051"),
  1040 => std_logic_vector'(x"81ff4002"),
  1041 => std_logic_vector'(x"610342b5"),
  1042 => std_logic_vector'(x"c164608c"),
  1043 => std_logic_vector'(x"c16c44f7"),
  1044 => std_logic_vector'(x"c16844f7"),
  1045 => std_logic_vector'(x"464d44f7"),
  1046 => std_logic_vector'(x"434a434a"),
  1047 => std_logic_vector'(x"443b434a"),
  1048 => std_logic_vector'(x"44f76011"),
  1049 => std_logic_vector'(x"44e8c168"),
  1050 => std_logic_vector'(x"60114009"),
  1051 => std_logic_vector'(x"c16c44f7"),
  1052 => std_logic_vector'(x"400944e8"),
  1053 => std_logic_vector'(x"c16444f7"),
  1054 => std_logic_vector'(x"608c04e8"),
  1055 => std_logic_vector'(x"c1646127"),
  1056 => std_logic_vector'(x"601144f7"),
  1057 => std_logic_vector'(x"28474007"),
  1058 => std_logic_vector'(x"005e6b1d"),
  1059 => std_logic_vector'(x"6011608c"),
  1060 => std_logic_vector'(x"62038002"),
  1061 => std_logic_vector'(x"620340d9"),
  1062 => std_logic_vector'(x"40934275"),
  1063 => std_logic_vector'(x"400d6b11"),
  1064 => std_logic_vector'(x"40932856"),
  1065 => std_logic_vector'(x"66008001"),
  1066 => std_logic_vector'(x"08416303"),
  1067 => std_logic_vector'(x"61036b1d"),
  1068 => std_logic_vector'(x"62038002"),
  1069 => std_logic_vector'(x"00e040d9"),
  1070 => std_logic_vector'(x"c9dc608c"),
  1071 => std_logic_vector'(x"ca28608c"),
  1072 => std_logic_vector'(x"ca54608c"),
  1073 => std_logic_vector'(x"ca68608c"),
  1074 => std_logic_vector'(x"8000608c"),
  1075 => std_logic_vector'(x"28694454"),
  1076 => std_logic_vector'(x"61270870"),
  1077 => std_logic_vector'(x"620340d9"),
  1078 => std_logic_vector'(x"44626b1d"),
  1079 => std_logic_vector'(x"08692870"),
  1080 => std_logic_vector'(x"479b43bc"),
  1081 => std_logic_vector'(x"608c0032"),
  1082 => std_logic_vector'(x"479bca88"),
  1083 => std_logic_vector'(x"6111c9dc"),
  1084 => std_logic_vector'(x"69038008"),
  1085 => std_logic_vector'(x"ca284865"),
  1086 => std_logic_vector'(x"80046111"),
  1087 => std_logic_vector'(x"80076903"),
  1088 => std_logic_vector'(x"48656303"),
  1089 => std_logic_vector'(x"6111ca54"),
  1090 => std_logic_vector'(x"69038002"),
  1091 => std_logic_vector'(x"63038003"),
  1092 => std_logic_vector'(x"ca684865"),
  1093 => std_logic_vector'(x"80036111"),
  1094 => std_logic_vector'(x"48656303"),
  1095 => std_logic_vector'(x"80804032"),
  1096 => std_logic_vector'(x"28946303"),
  1097 => std_logic_vector'(x"079bca8d"),
  1098 => std_logic_vector'(x"4113608c"),
  1099 => std_logic_vector'(x"608c0874"),
  1100 => std_logic_vector'(x"4028805a"),
  1101 => std_logic_vector'(x"074f4032"),
  1102 => std_logic_vector'(x"804a608c"),
  1103 => std_logic_vector'(x"40324028"),
  1104 => std_logic_vector'(x"608c074f"),
  1105 => std_logic_vector'(x"608cca9c"),
  1106 => std_logic_vector'(x"44f7c160"),
  1107 => std_logic_vector'(x"46134813"),
  1108 => std_logic_vector'(x"40dd8040"),
  1109 => std_logic_vector'(x"6011402e"),
  1110 => std_logic_vector'(x"6011474f"),
  1111 => std_logic_vector'(x"60114093"),
  1112 => std_logic_vector'(x"47558004"),
  1113 => std_logic_vector'(x"60114032"),
  1114 => std_logic_vector'(x"6903800f"),
  1115 => std_logic_vector'(x"ffff28c3"),
  1116 => std_logic_vector'(x"80246303"),
  1117 => std_logic_vector'(x"60114028"),
  1118 => std_logic_vector'(x"44e4474f"),
  1119 => std_logic_vector'(x"40288023"),
  1120 => std_logic_vector'(x"4813474f"),
  1121 => std_logic_vector'(x"601108cf"),
  1122 => std_logic_vector'(x"63039fff"),
  1123 => std_logic_vector'(x"61104111"),
  1124 => std_logic_vector'(x"6903800d"),
  1125 => std_logic_vector'(x"ca9c400b"),
  1126 => std_logic_vector'(x"44f76203"),
  1127 => std_logic_vector'(x"800242f8"),
  1128 => std_logic_vector'(x"40646203"),
  1129 => std_logic_vector'(x"28aa6703"),
  1130 => std_logic_vector'(x"c160405e"),
  1131 => std_logic_vector'(x"608c04e8"),
  1132 => std_logic_vector'(x"8000405e"),
  1133 => std_logic_vector'(x"012b608c"),
  1134 => std_logic_vector'(x"000b608c"),
  1135 => std_logic_vector'(x"40dd608c"),
  1136 => std_logic_vector'(x"28e34454"),
  1137 => std_logic_vector'(x"612708f7"),
  1138 => std_logic_vector'(x"408444ca"),
  1139 => std_logic_vector'(x"40846111"),
  1140 => std_logic_vector'(x"4060410a"),
  1141 => std_logic_vector'(x"401328f2"),
  1142 => std_logic_vector'(x"40024111"),
  1143 => std_logic_vector'(x"6b1d6003"),
  1144 => std_logic_vector'(x"608c43bc"),
  1145 => std_logic_vector'(x"6b1d4002"),
  1146 => std_logic_vector'(x"28f74462"),
  1147 => std_logic_vector'(x"43bc08e3"),
  1148 => std_logic_vector'(x"80006103"),
  1149 => std_logic_vector'(x"4053608c"),
  1150 => std_logic_vector'(x"61104064"),
  1151 => std_logic_vector'(x"6127410a"),
  1152 => std_logic_vector'(x"48df4078"),
  1153 => std_logic_vector'(x"29074060"),
  1154 => std_logic_vector'(x"61036b1d"),
  1155 => std_logic_vector'(x"6b1d608c"),
  1156 => std_logic_vector'(x"290d6011"),
  1157 => std_logic_vector'(x"41114011"),
  1158 => std_logic_vector'(x"608c0002"),
  1159 => std_logic_vector'(x"02cc8020"),
  1160 => std_logic_vector'(x"4064608c"),
  1161 => std_logic_vector'(x"40046203"),
  1162 => std_logic_vector'(x"80204084"),
  1163 => std_logic_vector'(x"61116703"),
  1164 => std_logic_vector'(x"291c6303"),
  1165 => std_logic_vector'(x"09114004"),
  1166 => std_logic_vector'(x"6011608c"),
  1167 => std_logic_vector'(x"29234007"),
  1168 => std_logic_vector'(x"0051405e"),
  1169 => std_logic_vector'(x"4638608c"),
  1170 => std_logic_vector'(x"60114064"),
  1171 => std_logic_vector'(x"4064293b"),
  1172 => std_logic_vector'(x"40534644"),
  1173 => std_logic_vector'(x"40786111"),
  1174 => std_logic_vector'(x"48fb4057"),
  1175 => std_logic_vector'(x"29384007"),
  1176 => std_logic_vector'(x"405e406d"),
  1177 => std_logic_vector'(x"6b1d6b1d"),
  1178 => std_logic_vector'(x"405e6110"),
  1179 => std_logic_vector'(x"608c0051"),
  1180 => std_logic_vector'(x"41248001"),
  1181 => std_logic_vector'(x"405e0925"),
  1182 => std_logic_vector'(x"6b1d6b1d"),
  1183 => std_logic_vector'(x"405e6110"),
  1184 => std_logic_vector'(x"608c8000"),
  1185 => std_logic_vector'(x"074f44f7"),
  1186 => std_logic_vector'(x"4121608c"),
  1187 => std_logic_vector'(x"6127294c"),
  1188 => std_logic_vector'(x"6b1d4945"),
  1189 => std_logic_vector'(x"074f6011"),
  1190 => std_logic_vector'(x"803c608c"),
  1191 => std_logic_vector'(x"41214028"),
  1192 => std_logic_vector'(x"47558000"),
  1193 => std_logic_vector'(x"4028803e"),
  1194 => std_logic_vector'(x"09454032"),
  1195 => std_logic_vector'(x"c160608c"),
  1196 => std_logic_vector'(x"611044f7"),
  1197 => std_logic_vector'(x"414a4813"),
  1198 => std_logic_vector'(x"471c470b"),
  1199 => std_logic_vector'(x"4735471c"),
  1200 => std_logic_vector'(x"403240e0"),
  1201 => std_logic_vector'(x"04e8c160"),
  1202 => std_logic_vector'(x"4060608c"),
  1203 => std_logic_vector'(x"c16029a6"),
  1204 => std_logic_vector'(x"612744f7"),
  1205 => std_logic_vector'(x"40044813"),
  1206 => std_logic_vector'(x"69038004"),
  1207 => std_logic_vector'(x"80004002"),
  1208 => std_logic_vector'(x"61274448"),
  1209 => std_logic_vector'(x"6011402e"),
  1210 => std_logic_vector'(x"80086011"),
  1211 => std_logic_vector'(x"4032475a"),
  1212 => std_logic_vector'(x"80104032"),
  1213 => std_logic_vector'(x"44488000"),
  1214 => std_logic_vector'(x"60116127"),
  1215 => std_logic_vector'(x"49574084"),
  1216 => std_logic_vector'(x"6b1d4002"),
  1217 => std_logic_vector'(x"29854462"),
  1218 => std_logic_vector'(x"43bc097c"),
  1219 => std_logic_vector'(x"61104032"),
  1220 => std_logic_vector'(x"80008010"),
  1221 => std_logic_vector'(x"61274448"),
  1222 => std_logic_vector'(x"40846011"),
  1223 => std_logic_vector'(x"80206011"),
  1224 => std_logic_vector'(x"47d2807f"),
  1225 => std_logic_vector'(x"29966600"),
  1226 => std_logic_vector'(x"802e6103"),
  1227 => std_logic_vector'(x"40024028"),
  1228 => std_logic_vector'(x"44626b1d"),
  1229 => std_logic_vector'(x"098b299c"),
  1230 => std_logic_vector'(x"610343bc"),
  1231 => std_logic_vector'(x"44626b1d"),
  1232 => std_logic_vector'(x"097129a2"),
  1233 => std_logic_vector'(x"6b1d43bc"),
  1234 => std_logic_vector'(x"44e8c160"),
  1235 => std_logic_vector'(x"608c6103"),
  1236 => std_logic_vector'(x"43118001"),
  1237 => std_logic_vector'(x"29cc6011"),
  1238 => std_logic_vector'(x"cb524064"),
  1239 => std_logic_vector'(x"48fb40d9"),
  1240 => std_logic_vector'(x"29b54007"),
  1241 => std_logic_vector'(x"4002405e"),
  1242 => std_logic_vector'(x"406409c7"),
  1243 => std_logic_vector'(x"40d9cb57"),
  1244 => std_logic_vector'(x"400748fb"),
  1245 => std_logic_vector'(x"405e29c1"),
  1246 => std_logic_vector'(x"60114004"),
  1247 => std_logic_vector'(x"400229c0"),
  1248 => std_logic_vector'(x"cb5e09c7"),
  1249 => std_logic_vector'(x"48fb40d9"),
  1250 => std_logic_vector'(x"29c74007"),
  1251 => std_logic_vector'(x"40604004"),
  1252 => std_logic_vector'(x"29cb4007"),
  1253 => std_logic_vector'(x"09a9608c"),
  1254 => std_logic_vector'(x"45c4405e"),
  1255 => std_logic_vector'(x"29a94007"),
  1256 => std_logic_vector'(x"608c6103"),
  1257 => std_logic_vector'(x"29d54007"),
  1258 => std_logic_vector'(x"608c09a8"),
  1259 => std_logic_vector'(x"07c4608c"),
  1260 => std_logic_vector'(x"07bb608c"),
  1261 => std_logic_vector'(x"4311608c"),
  1262 => std_logic_vector'(x"6003428b"),
  1263 => std_logic_vector'(x"40604015"),
  1264 => std_logic_vector'(x"608c6303"),
  1265 => std_logic_vector'(x"000749db"),
  1266 => std_logic_vector'(x"464d608c"),
  1267 => std_logic_vector'(x"434a89d0"),
  1268 => std_logic_vector'(x"443b434a"),
  1269 => std_logic_vector'(x"04f74009"),
  1270 => std_logic_vector'(x"464d608c"),
  1271 => std_logic_vector'(x"434a82a6"),
  1272 => std_logic_vector'(x"434a434a"),
  1273 => std_logic_vector'(x"4009443b"),
  1274 => std_logic_vector'(x"608c014c"),
  1275 => std_logic_vector'(x"46534613"),
  1276 => std_logic_vector'(x"40096011"),
  1277 => std_logic_vector'(x"44f7c18c"),
  1278 => std_logic_vector'(x"45242a01"),
  1279 => std_logic_vector'(x"442344f7"),
  1280 => std_logic_vector'(x"61100a04"),
  1281 => std_logic_vector'(x"02f844f7"),
  1282 => std_logic_vector'(x"cbe0608c"),
  1283 => std_logic_vector'(x"6110608c"),
  1284 => std_logic_vector'(x"cbe02a0f"),
  1285 => std_logic_vector'(x"800144e8"),
  1286 => std_logic_vector'(x"450c6600"),
  1287 => std_logic_vector'(x"61030a10"),
  1288 => std_logic_vector'(x"478f608c"),
  1289 => std_logic_vector'(x"0423940e"),
  1290 => std_logic_vector'(x"801b608c"),
  1291 => std_logic_vector'(x"805b4028"),
  1292 => std_logic_vector'(x"608c0028"),
  1293 => std_logic_vector'(x"40024a15"),
  1294 => std_logic_vector'(x"475a8000"),
  1295 => std_logic_vector'(x"4028803b"),
  1296 => std_logic_vector'(x"80004002"),
  1297 => std_logic_vector'(x"8048475a"),
  1298 => std_logic_vector'(x"608c0028"),
  1299 => std_logic_vector'(x"80008000"),
  1300 => std_logic_vector'(x"4a154a1a"),
  1301 => std_logic_vector'(x"0028804a"),
  1302 => std_logic_vector'(x"608c608c"),
  1303 => std_logic_vector'(x"608c608c"),
  1304 => std_logic_vector'(x"4084405c"),
  1305 => std_logic_vector'(x"61106203"),
  1306 => std_logic_vector'(x"608c00c4"),
  1307 => std_logic_vector'(x"40d9405c"),
  1308 => std_logic_vector'(x"40c46203"),
  1309 => std_logic_vector'(x"61108001"),
  1310 => std_logic_vector'(x"608c0a30"),
  1311 => std_logic_vector'(x"405c6127"),
  1312 => std_logic_vector'(x"40d96b11"),
  1313 => std_logic_vector'(x"61106203"),
  1314 => std_logic_vector'(x"6b1d42d8"),
  1315 => std_logic_vector'(x"608c0a30"),
  1316 => std_logic_vector'(x"44f7c160"),
  1317 => std_logic_vector'(x"48136127"),
  1318 => std_logic_vector'(x"80008000"),
  1319 => std_logic_vector'(x"61034072"),
  1320 => std_logic_vector'(x"42b58002"),
  1321 => std_logic_vector'(x"6103405e"),
  1322 => std_logic_vector'(x"80026127"),
  1323 => std_logic_vector'(x"6b1d4124"),
  1324 => std_logic_vector'(x"c1606b1d"),
  1325 => std_logic_vector'(x"608c04e8"),
  1326 => std_logic_vector'(x"608ccc88"),
  1327 => std_logic_vector'(x"608cccac"),
  1328 => std_logic_vector'(x"40076111"),
  1329 => std_logic_vector'(x"61032a65"),
  1330 => std_logic_vector'(x"6127608c"),
  1331 => std_logic_vector'(x"40846111"),
  1332 => std_logic_vector'(x"67038078"),
  1333 => std_logic_vector'(x"80012a71"),
  1334 => std_logic_vector'(x"4a484124"),
  1335 => std_logic_vector'(x"0a366b1d"),
  1336 => std_logic_vector'(x"6111608c"),
  1337 => std_logic_vector'(x"806d4084"),
  1338 => std_logic_vector'(x"2a7f6703"),
  1339 => std_logic_vector'(x"41248001"),
  1340 => std_logic_vector'(x"6b11800d"),
  1341 => std_logic_vector'(x"800a4a36"),
  1342 => std_logic_vector'(x"0a366b1d"),
  1343 => std_logic_vector'(x"6111608c"),
  1344 => std_logic_vector'(x"806e4084"),
  1345 => std_logic_vector'(x"2a8b6703"),
  1346 => std_logic_vector'(x"41248001"),
  1347 => std_logic_vector'(x"40d9ccac"),
  1348 => std_logic_vector'(x"0a3e6b1d"),
  1349 => std_logic_vector'(x"6111608c"),
  1350 => std_logic_vector'(x"80614084"),
  1351 => std_logic_vector'(x"4002807a"),
  1352 => std_logic_vector'(x"2a9c47d2"),
  1353 => std_logic_vector'(x"40846111"),
  1354 => std_logic_vector'(x"410a8061"),
  1355 => std_logic_vector'(x"6203cc88"),
  1356 => std_logic_vector'(x"6b1d4084"),
  1357 => std_logic_vector'(x"0aa04a36"),
  1358 => std_logic_vector'(x"40846111"),
  1359 => std_logic_vector'(x"4a366b1d"),
  1360 => std_logic_vector'(x"01248001"),
  1361 => std_logic_vector'(x"6011608c"),
  1362 => std_logic_vector'(x"80006127"),
  1363 => std_logic_vector'(x"40c46110"),
  1364 => std_logic_vector'(x"2ac06011"),
  1365 => std_logic_vector'(x"40846111"),
  1366 => std_logic_vector'(x"400d8022"),
  1367 => std_logic_vector'(x"61112ac0"),
  1368 => std_logic_vector'(x"805c4084"),
  1369 => std_logic_vector'(x"2ab96703"),
  1370 => std_logic_vector'(x"41248001"),
  1371 => std_logic_vector'(x"4a606b11"),
  1372 => std_logic_vector'(x"61110abf"),
  1373 => std_logic_vector'(x"6b114084"),
  1374 => std_logic_vector'(x"80014a36"),
  1375 => std_logic_vector'(x"0aa84124"),
  1376 => std_logic_vector'(x"2ac46011"),
  1377 => std_logic_vector'(x"41248001"),
  1378 => std_logic_vector'(x"61036b1d"),
  1379 => std_logic_vector'(x"42fa608c"),
  1380 => std_logic_vector'(x"44f7c188"),
  1381 => std_logic_vector'(x"405c4124"),
  1382 => std_logic_vector'(x"4aa3c908"),
  1383 => std_logic_vector'(x"410a6003"),
  1384 => std_logic_vector'(x"4066c188"),
  1385 => std_logic_vector'(x"608cc908"),
  1386 => std_logic_vector'(x"40d94ac7"),
  1387 => std_logic_vector'(x"44f7c18c"),
  1388 => std_logic_vector'(x"07952ada"),
  1389 => std_logic_vector'(x"464d608c"),
  1390 => std_logic_vector'(x"434a8c1e"),
  1391 => std_logic_vector'(x"44f7443b"),
  1392 => std_logic_vector'(x"608c02f8"),
  1393 => std_logic_vector'(x"04f74653"),
  1394 => std_logic_vector'(x"4653608c"),
  1395 => std_logic_vector'(x"608c04e8"),
  1396 => std_logic_vector'(x"44f7c18c"),
  1397 => std_logic_vector'(x"461b2aef"),
  1398 => std_logic_vector'(x"442395ca"),
  1399 => std_logic_vector'(x"46130af1"),
  1400 => std_logic_vector'(x"608c0ae5"),
  1401 => std_logic_vector'(x"44f7c18c"),
  1402 => std_logic_vector'(x"461b2af9"),
  1403 => std_logic_vector'(x"442395c4"),
  1404 => std_logic_vector'(x"46130afb"),
  1405 => std_logic_vector'(x"608c0ae2"),
  1406 => std_logic_vector'(x"2b046011"),
  1407 => std_logic_vector'(x"40644004"),
  1408 => std_logic_vector'(x"40846203"),
  1409 => std_logic_vector'(x"0afc470f"),
  1410 => std_logic_vector'(x"608c005e"),
  1411 => std_logic_vector'(x"0348464d"),
  1412 => std_logic_vector'(x"464d608c"),
  1413 => std_logic_vector'(x"8000411e"),
  1414 => std_logic_vector'(x"434a8000"),
  1415 => std_logic_vector'(x"04f7443b"),
  1416 => std_logic_vector'(x"6110608c"),
  1417 => std_logic_vector'(x"608c04e8"),
  1418 => std_logic_vector'(x"6111464d"),
  1419 => std_logic_vector'(x"6203434a"),
  1420 => std_logic_vector'(x"44f7443b"),
  1421 => std_logic_vector'(x"608c6203"),
  1422 => std_logic_vector'(x"60008001"),
  1423 => std_logic_vector'(x"608c0b14"),
  1424 => std_logic_vector'(x"8001412b"),
  1425 => std_logic_vector'(x"0b14400b"),
  1426 => std_logic_vector'(x"48db608c"),
  1427 => std_logic_vector'(x"48dd8001"),
  1428 => std_logic_vector'(x"608c0b14"),
  1429 => std_logic_vector'(x"8000608c"),
  1430 => std_logic_vector'(x"04e86110"),
  1431 => std_logic_vector'(x"4051608c"),
  1432 => std_logic_vector'(x"04e86110"),
  1433 => std_logic_vector'(x"cdac608c"),
  1434 => std_logic_vector'(x"6011608c"),
  1435 => std_logic_vector'(x"64034007"),
  1436 => std_logic_vector'(x"04e8cdac"),
  1437 => std_logic_vector'(x"cdac608c"),
  1438 => std_logic_vector'(x"601144f7"),
  1439 => std_logic_vector'(x"6a03800d"),
  1440 => std_logic_vector'(x"60116503"),
  1441 => std_logic_vector'(x"69038011"),
  1442 => std_logic_vector'(x"60116503"),
  1443 => std_logic_vector'(x"6a038005"),
  1444 => std_logic_vector'(x"60116503"),
  1445 => std_logic_vector'(x"04e8cdac"),
  1446 => std_logic_vector'(x"4b3b608c"),
  1447 => std_logic_vector'(x"600341aa"),
  1448 => std_logic_vector'(x"0007608c"),
  1449 => std_logic_vector'(x"464d608c"),
  1450 => std_logic_vector'(x"434a6111"),
  1451 => std_logic_vector'(x"40096110"),
  1452 => std_logic_vector'(x"443b6110"),
  1453 => std_logic_vector'(x"611144f7"),
  1454 => std_logic_vector'(x"620344f7"),
  1455 => std_logic_vector'(x"02f844f7"),
  1456 => std_logic_vector'(x"464d608c"),
  1457 => std_logic_vector'(x"434a6111"),
  1458 => std_logic_vector'(x"443b6203"),
  1459 => std_logic_vector'(x"620344f7"),
  1460 => std_logic_vector'(x"6011608c"),
  1461 => std_logic_vector'(x"608c014c"),
  1462 => std_logic_vector'(x"411e464d"),
  1463 => std_logic_vector'(x"434a6127"),
  1464 => std_logic_vector'(x"434a6011"),
  1465 => std_logic_vector'(x"400b8002"),
  1466 => std_logic_vector'(x"2b774454"),
  1467 => std_logic_vector'(x"61270b7f"),
  1468 => std_logic_vector'(x"434a9654"),
  1469 => std_logic_vector'(x"400b8001"),
  1470 => std_logic_vector'(x"44906b1d"),
  1471 => std_logic_vector'(x"43bc2b77"),
  1472 => std_logic_vector'(x"60114009"),
  1473 => std_logic_vector'(x"6b1d4009"),
  1474 => std_logic_vector'(x"44f74053"),
  1475 => std_logic_vector'(x"400b8002"),
  1476 => std_logic_vector'(x"075e4124"),
  1477 => std_logic_vector'(x"4613608c"),
  1478 => std_logic_vector'(x"44f74653"),
  1479 => std_logic_vector'(x"608c6203"),
  1480 => std_logic_vector'(x"04f74b8b"),
  1481 => std_logic_vector'(x"4b8b608c"),
  1482 => std_logic_vector'(x"608c04e8"),
  1483 => std_logic_vector'(x"411e4633"),
  1484 => std_logic_vector'(x"44f76111"),
  1485 => std_logic_vector'(x"405c4348"),
  1486 => std_logic_vector'(x"608c04e8"),
  1487 => std_logic_vector'(x"04234b90"),
  1488 => std_logic_vector'(x"ce48608c"),
  1489 => std_logic_vector'(x"8000608c"),
  1490 => std_logic_vector'(x"8001608c"),
  1491 => std_logic_vector'(x"8100608c"),
  1492 => std_logic_vector'(x"04f96203"),
  1493 => std_logic_vector'(x"04fb608c"),
  1494 => std_logic_vector'(x"04f9608c"),
  1495 => std_logic_vector'(x"8001608c"),
  1496 => std_logic_vector'(x"4ba76111"),
  1497 => std_logic_vector'(x"61118000"),
  1498 => std_logic_vector'(x"800144f9"),
  1499 => std_logic_vector'(x"44f96111"),
  1500 => std_logic_vector'(x"608c0bb2"),
  1501 => std_logic_vector'(x"61108000"),
  1502 => std_logic_vector'(x"608c04f9"),
  1503 => std_logic_vector'(x"61108001"),
  1504 => std_logic_vector'(x"608c04f9"),
  1505 => std_logic_vector'(x"608c800b"),
  1506 => std_logic_vector'(x"608c800c"),
  1507 => std_logic_vector'(x"608c800d"),
  1508 => std_logic_vector'(x"800b6903"),
  1509 => std_logic_vector'(x"800144f9"),
  1510 => std_logic_vector'(x"44f9800d"),
  1511 => std_logic_vector'(x"800d8000"),
  1512 => std_logic_vector'(x"608c04f9"),
  1513 => std_logic_vector'(x"80088000"),
  1514 => std_logic_vector'(x"44488000"),
  1515 => std_logic_vector'(x"61116127"),
  1516 => std_logic_vector'(x"69038007"),
  1517 => std_logic_vector'(x"44f9800b"),
  1518 => std_logic_vector'(x"4bbe800d"),
  1519 => std_logic_vector'(x"800c4111"),
  1520 => std_logic_vector'(x"620344fb"),
  1521 => std_logic_vector'(x"4bba800d"),
  1522 => std_logic_vector'(x"41116110"),
  1523 => std_logic_vector'(x"6b1d6110"),
  1524 => std_logic_vector'(x"2beb4462"),
  1525 => std_logic_vector'(x"43bc0bd6"),
  1526 => std_logic_vector'(x"608c6003"),
  1527 => std_logic_vector'(x"0bd28000"),
  1528 => std_logic_vector'(x"8001608c"),
  1529 => std_logic_vector'(x"4ba7800b"),
  1530 => std_logic_vector'(x"800d8001"),
  1531 => std_logic_vector'(x"608c0ba7"),
  1532 => std_logic_vector'(x"80076011"),
  1533 => std_logic_vector'(x"60114bc8"),
  1534 => std_logic_vector'(x"4bc88006"),
  1535 => std_logic_vector'(x"80056011"),
  1536 => std_logic_vector'(x"60114bc8"),
  1537 => std_logic_vector'(x"4bc88004"),
  1538 => std_logic_vector'(x"80036011"),
  1539 => std_logic_vector'(x"60114bc8"),
  1540 => std_logic_vector'(x"4bc88002"),
  1541 => std_logic_vector'(x"80016011"),
  1542 => std_logic_vector'(x"80004bc8"),
  1543 => std_logic_vector'(x"608c0bc8"),
  1544 => std_logic_vector'(x"444840dd"),
  1545 => std_logic_vector'(x"44ca6127"),
  1546 => std_logic_vector'(x"4bf84084"),
  1547 => std_logic_vector'(x"44626b1d"),
  1548 => std_logic_vector'(x"0c122c1a"),
  1549 => std_logic_vector'(x"608c43bc"),
  1550 => std_logic_vector'(x"04fb9010"),
  1551 => std_logic_vector'(x"8000608c"),
  1552 => std_logic_vector'(x"44f99010"),
  1553 => std_logic_vector'(x"44fb9014"),
  1554 => std_logic_vector'(x"04fb9018"),
  1555 => std_logic_vector'(x"4c1f608c"),
  1556 => std_logic_vector'(x"4c1c4053"),
  1557 => std_logic_vector'(x"608c06b5"),
  1558 => std_logic_vector'(x"04fb901c"),
  1559 => std_logic_vector'(x"801e608c"),
  1560 => std_logic_vector'(x"6a03800f"),
  1561 => std_logic_vector'(x"6403c240"),
  1562 => std_logic_vector'(x"608c0c27"),
  1563 => std_logic_vector'(x"800ff735"),
  1564 => std_logic_vector'(x"ca006a03"),
  1565 => std_logic_vector'(x"0c276403"),
  1566 => std_logic_vector'(x"414a608c"),
  1567 => std_logic_vector'(x"83e84c1c"),
  1568 => std_logic_vector'(x"4c1f46b5"),
  1569 => std_logic_vector'(x"40644130"),
  1570 => std_logic_vector'(x"41674c1f"),
  1571 => std_logic_vector'(x"005e2c43"),
  1572 => std_logic_vector'(x"cf50608c"),
  1573 => std_logic_vector'(x"05d240d9"),
  1574 => std_logic_vector'(x"cf64608c"),
  1575 => std_logic_vector'(x"cf7c0830"),
  1576 => std_logic_vector'(x"8001608c"),
  1577 => std_logic_vector'(x"6a03800f"),
  1578 => std_logic_vector'(x"6403ffff"),
  1579 => std_logic_vector'(x"6a03800f"),
  1580 => std_logic_vector'(x"6403ffff"),
  1581 => std_logic_vector'(x"608c6600"),
  1582 => std_logic_vector'(x"61114053"),
  1583 => std_logic_vector'(x"67036111"),
  1584 => std_logic_vector'(x"61032c65"),
  1585 => std_logic_vector'(x"6f036103"),
  1586 => std_logic_vector'(x"40170c6a"),
  1587 => std_logic_vector'(x"61036127"),
  1588 => std_logic_vector'(x"6b1d6103"),
  1589 => std_logic_vector'(x"8000608c"),
  1590 => std_logic_vector'(x"80006110"),
  1591 => std_logic_vector'(x"61274448"),
  1592 => std_logic_vector'(x"61116103"),
  1593 => std_logic_vector'(x"611144f7"),
  1594 => std_logic_vector'(x"401744f7"),
  1595 => std_logic_vector'(x"80002c7a"),
  1596 => std_logic_vector'(x"0c906b1d"),
  1597 => std_logic_vector'(x"44f76111"),
  1598 => std_logic_vector'(x"44f76111"),
  1599 => std_logic_vector'(x"60116f03"),
  1600 => std_logic_vector'(x"6b1d2c83"),
  1601 => std_logic_vector'(x"40530c90"),
  1602 => std_logic_vector'(x"400b8001"),
  1603 => std_logic_vector'(x"40536203"),
  1604 => std_logic_vector'(x"400b8001"),
  1605 => std_logic_vector'(x"40536203"),
  1606 => std_logic_vector'(x"44626b1d"),
  1607 => std_logic_vector'(x"0c6f2c90"),
  1608 => std_logic_vector'(x"405743bc"),
  1609 => std_logic_vector'(x"608c005e"),
  1610 => std_logic_vector'(x"61116110"),
  1611 => std_logic_vector'(x"400b4004"),
  1612 => std_logic_vector'(x"40576203"),
  1613 => std_logic_vector'(x"61116110"),
  1614 => std_logic_vector'(x"400b4004"),
  1615 => std_logic_vector'(x"40576203"),
  1616 => std_logic_vector'(x"61108001"),
  1617 => std_logic_vector'(x"44488000"),
  1618 => std_logic_vector'(x"61116127"),
  1619 => std_logic_vector'(x"800044f7"),
  1620 => std_logic_vector'(x"65036600"),
  1621 => std_logic_vector'(x"40538000"),
  1622 => std_logic_vector'(x"41308000"),
  1623 => std_logic_vector'(x"47c48003"),
  1624 => std_logic_vector'(x"800044f7"),
  1625 => std_logic_vector'(x"61104130"),
  1626 => std_logic_vector'(x"47c48003"),
  1627 => std_logic_vector'(x"405344e8"),
  1628 => std_logic_vector'(x"400b8001"),
  1629 => std_logic_vector'(x"4053410a"),
  1630 => std_logic_vector'(x"400b8001"),
  1631 => std_logic_vector'(x"4053410a"),
  1632 => std_logic_vector'(x"44626b1d"),
  1633 => std_logic_vector'(x"0ca42cc4"),
  1634 => std_logic_vector'(x"610343bc"),
  1635 => std_logic_vector'(x"608c005e"),
  1636 => std_logic_vector'(x"40578000"),
  1637 => std_logic_vector'(x"44488000"),
  1638 => std_logic_vector'(x"60116127"),
  1639 => std_logic_vector'(x"601144f7"),
  1640 => std_logic_vector'(x"80016127"),
  1641 => std_logic_vector'(x"40536903"),
  1642 => std_logic_vector'(x"61116403"),
  1643 => std_logic_vector'(x"400944e8"),
  1644 => std_logic_vector'(x"80016b1d"),
  1645 => std_logic_vector'(x"41086303"),
  1646 => std_logic_vector'(x"80016011"),
  1647 => std_logic_vector'(x"65036903"),
  1648 => std_logic_vector'(x"6b1d6110"),
  1649 => std_logic_vector'(x"2ce54462"),
  1650 => std_logic_vector'(x"43bc0ccc"),
  1651 => std_logic_vector'(x"61036103"),
  1652 => std_logic_vector'(x"8000608c"),
  1653 => std_logic_vector'(x"40648000"),
  1654 => std_logic_vector'(x"4153cf7c"),
  1655 => std_logic_vector'(x"8002cf7c"),
  1656 => std_logic_vector'(x"6203400b"),
  1657 => std_logic_vector'(x"61274153"),
  1658 => std_logic_vector'(x"61106127"),
  1659 => std_logic_vector'(x"6b116011"),
  1660 => std_logic_vector'(x"cf7c41aa"),
  1661 => std_logic_vector'(x"400b8002"),
  1662 => std_logic_vector'(x"41536203"),
  1663 => std_logic_vector'(x"6b1d6111"),
  1664 => std_logic_vector'(x"cf7c41aa"),
  1665 => std_logic_vector'(x"400b8001"),
  1666 => std_logic_vector'(x"414c6203"),
  1667 => std_logic_vector'(x"cf7c4130"),
  1668 => std_logic_vector'(x"400b8001"),
  1669 => std_logic_vector'(x"41536203"),
  1670 => std_logic_vector'(x"41aa6b11"),
  1671 => std_logic_vector'(x"46444638"),
  1672 => std_logic_vector'(x"8001cf7c"),
  1673 => std_logic_vector'(x"6203400b"),
  1674 => std_logic_vector'(x"4130414c"),
  1675 => std_logic_vector'(x"cf7c4064"),
  1676 => std_logic_vector'(x"400b8001"),
  1677 => std_logic_vector'(x"41536203"),
  1678 => std_logic_vector'(x"6b1d6b1d"),
  1679 => std_logic_vector'(x"4c5c6110"),
  1680 => std_logic_vector'(x"cf7c2d26"),
  1681 => std_logic_vector'(x"400244f7"),
  1682 => std_logic_vector'(x"44e8cf7c"),
  1683 => std_logic_vector'(x"41aa6b1d"),
  1684 => std_logic_vector'(x"414ccf7c"),
  1685 => std_logic_vector'(x"cf7c4130"),
  1686 => std_logic_vector'(x"608c0153"),
  1687 => std_logic_vector'(x"608ccfcc"),
  1688 => std_logic_vector'(x"479bcfe8"),
  1689 => std_logic_vector'(x"6011cfcc"),
  1690 => std_logic_vector'(x"475244f7"),
  1691 => std_logic_vector'(x"60114009"),
  1692 => std_logic_vector'(x"475244f7"),
  1693 => std_logic_vector'(x"60114009"),
  1694 => std_logic_vector'(x"475244f7"),
  1695 => std_logic_vector'(x"44f74009"),
  1696 => std_logic_vector'(x"002e4752"),
  1697 => std_logic_vector'(x"cffc608c"),
  1698 => std_logic_vector'(x"cf7c479b"),
  1699 => std_logic_vector'(x"44f76011"),
  1700 => std_logic_vector'(x"40094752"),
  1701 => std_logic_vector'(x"44f76011"),
  1702 => std_logic_vector'(x"40094752"),
  1703 => std_logic_vector'(x"44f76011"),
  1704 => std_logic_vector'(x"40094752"),
  1705 => std_logic_vector'(x"475244f7"),
  1706 => std_logic_vector'(x"608c002e"),
  1707 => std_logic_vector'(x"cf7c4064"),
  1708 => std_logic_vector'(x"406d414c"),
  1709 => std_logic_vector'(x"2d824c5c"),
  1710 => std_logic_vector'(x"4153cfcc"),
  1711 => std_logic_vector'(x"80008000"),
  1712 => std_logic_vector'(x"8002cfcc"),
  1713 => std_logic_vector'(x"6203400b"),
  1714 => std_logic_vector'(x"80004153"),
  1715 => std_logic_vector'(x"80408000"),
  1716 => std_logic_vector'(x"44488000"),
  1717 => std_logic_vector'(x"41836127"),
  1718 => std_logic_vector'(x"8004cfcc"),
  1719 => std_logic_vector'(x"cfcc4cc8"),
  1720 => std_logic_vector'(x"8004cf7c"),
  1721 => std_logic_vector'(x"2d7c4c6b"),
  1722 => std_logic_vector'(x"40538001"),
  1723 => std_logic_vector'(x"61106403"),
  1724 => std_logic_vector'(x"cfcccf7c"),
  1725 => std_logic_vector'(x"4c948004"),
  1726 => std_logic_vector'(x"44626b1d"),
  1727 => std_logic_vector'(x"0d6a2d80"),
  1728 => std_logic_vector'(x"0d8643bc"),
  1729 => std_logic_vector'(x"479bd00c"),
  1730 => std_logic_vector'(x"050c8088"),
  1731 => std_logic_vector'(x"cf7c608c"),
  1732 => std_logic_vector'(x"6110414c"),
  1733 => std_logic_vector'(x"8002cf7c"),
  1734 => std_logic_vector'(x"6203400b"),
  1735 => std_logic_vector'(x"6110414c"),
  1736 => std_logic_vector'(x"e100608c"),
  1737 => std_logic_vector'(x"6011608c"),
  1738 => std_logic_vector'(x"050c474f"),
  1739 => std_logic_vector'(x"80c8608c"),
  1740 => std_logic_vector'(x"44f9e100"),
  1741 => std_logic_vector'(x"e1008000"),
  1742 => std_logic_vector'(x"62038001"),
  1743 => std_logic_vector'(x"808044f9"),
  1744 => std_logic_vector'(x"8002e100"),
  1745 => std_logic_vector'(x"04f96203"),
  1746 => std_logic_vector'(x"e100608c"),
  1747 => std_logic_vector'(x"62038003"),
  1748 => std_logic_vector'(x"808044f9"),
  1749 => std_logic_vector'(x"64038010"),
  1750 => std_logic_vector'(x"8004e100"),
  1751 => std_logic_vector'(x"44f96203"),
  1752 => std_logic_vector'(x"8004e100"),
  1753 => std_logic_vector'(x"44fb6203"),
  1754 => std_logic_vector'(x"80026011"),
  1755 => std_logic_vector'(x"2dba6303"),
  1756 => std_logic_vector'(x"0db06103"),
  1757 => std_logic_vector'(x"63038080"),
  1758 => std_logic_vector'(x"80852dbf"),
  1759 => std_logic_vector'(x"608c0d93"),
  1760 => std_logic_vector'(x"4da54111"),
  1761 => std_logic_vector'(x"8003e100"),
  1762 => std_logic_vector'(x"44f96203"),
  1763 => std_logic_vector'(x"80108040"),
  1764 => std_logic_vector'(x"e1006403"),
  1765 => std_logic_vector'(x"62038004"),
  1766 => std_logic_vector'(x"e10044f9"),
  1767 => std_logic_vector'(x"62038004"),
  1768 => std_logic_vector'(x"601144fb"),
  1769 => std_logic_vector'(x"63038002"),
  1770 => std_logic_vector'(x"61032dd7"),
  1771 => std_logic_vector'(x"80800dcd"),
  1772 => std_logic_vector'(x"2ddc6303"),
  1773 => std_logic_vector'(x"0d938086"),
  1774 => std_logic_vector'(x"4111608c"),
  1775 => std_logic_vector'(x"4da54002"),
  1776 => std_logic_vector'(x"80208040"),
  1777 => std_logic_vector'(x"80086403"),
  1778 => std_logic_vector'(x"e1006403"),
  1779 => std_logic_vector'(x"62038004"),
  1780 => std_logic_vector'(x"e10044f9"),
  1781 => std_logic_vector'(x"62038004"),
  1782 => std_logic_vector'(x"601144fb"),
  1783 => std_logic_vector'(x"63038002"),
  1784 => std_logic_vector'(x"61032df3"),
  1785 => std_logic_vector'(x"61030de9"),
  1786 => std_logic_vector'(x"8003e100"),
  1787 => std_logic_vector'(x"04fb6203"),
  1788 => std_logic_vector'(x"4111608c"),
  1789 => std_logic_vector'(x"60114da5"),
  1790 => std_logic_vector'(x"61104084"),
  1791 => std_logic_vector'(x"61104002"),
  1792 => std_logic_vector'(x"2e246011"),
  1793 => std_logic_vector'(x"40846111"),
  1794 => std_logic_vector'(x"8003e100"),
  1795 => std_logic_vector'(x"44f96203"),
  1796 => std_logic_vector'(x"60114004"),
  1797 => std_logic_vector'(x"80102e0d"),
  1798 => std_logic_vector'(x"80400e10"),
  1799 => std_logic_vector'(x"64038010"),
  1800 => std_logic_vector'(x"8004e100"),
  1801 => std_logic_vector'(x"44f96203"),
  1802 => std_logic_vector'(x"8004e100"),
  1803 => std_logic_vector'(x"44fb6203"),
  1804 => std_logic_vector'(x"80026011"),
  1805 => std_logic_vector'(x"2e1e6303"),
  1806 => std_logic_vector'(x"0e146103"),
  1807 => std_logic_vector'(x"63038080"),
  1808 => std_logic_vector'(x"80862e23"),
  1809 => std_logic_vector'(x"0dfd4d93"),
  1810 => std_logic_vector'(x"608c005e"),
  1811 => std_logic_vector'(x"40024111"),
  1812 => std_logic_vector'(x"60114da5"),
  1813 => std_logic_vector'(x"80014002"),
  1814 => std_logic_vector'(x"61274448"),
  1815 => std_logic_vector'(x"44ca6011"),
  1816 => std_logic_vector'(x"2e386703"),
  1817 => std_logic_vector'(x"80208040"),
  1818 => std_logic_vector'(x"80086403"),
  1819 => std_logic_vector'(x"0e396403"),
  1820 => std_logic_vector'(x"e1008020"),
  1821 => std_logic_vector'(x"62038004"),
  1822 => std_logic_vector'(x"e10044f9"),
  1823 => std_logic_vector'(x"62038004"),
  1824 => std_logic_vector'(x"601144fb"),
  1825 => std_logic_vector'(x"63038002"),
  1826 => std_logic_vector'(x"61032e47"),
  1827 => std_logic_vector'(x"40530e3d"),
  1828 => std_logic_vector'(x"611144ca"),
  1829 => std_logic_vector'(x"601140c4"),
  1830 => std_logic_vector'(x"620344ca"),
  1831 => std_logic_vector'(x"8003e100"),
  1832 => std_logic_vector'(x"44fb6203"),
  1833 => std_logic_vector'(x"40c46110"),
  1834 => std_logic_vector'(x"80804057"),
  1835 => std_logic_vector'(x"2e5a6303"),
  1836 => std_logic_vector'(x"0e5e6b1d"),
  1837 => std_logic_vector'(x"44626b1d"),
  1838 => std_logic_vector'(x"0e2d2e5e"),
  1839 => std_logic_vector'(x"610343bc"),
  1840 => std_logic_vector'(x"608c6103"),
  1841 => std_logic_vector'(x"608c8100"),
  1842 => std_logic_vector'(x"608c8101"),
  1843 => std_logic_vector'(x"608c8102"),
  1844 => std_logic_vector'(x"608c8180"),
  1845 => std_logic_vector'(x"608c8181"),
  1846 => std_logic_vector'(x"608c8182"),
  1847 => std_logic_vector'(x"608c8183"),
  1848 => std_logic_vector'(x"608c8190"),
  1849 => std_logic_vector'(x"608c8191"),
  1850 => std_logic_vector'(x"608c8192"),
  1851 => std_logic_vector'(x"608c8193"),
  1852 => std_logic_vector'(x"608c8201"),
  1853 => std_logic_vector'(x"04f98201"),
  1854 => std_logic_vector'(x"8070608c"),
  1855 => std_logic_vector'(x"800a608c"),
  1856 => std_logic_vector'(x"800c608c"),
  1857 => std_logic_vector'(x"d17c608c"),
  1858 => std_logic_vector'(x"6011608c"),
  1859 => std_logic_vector'(x"4dc04057"),
  1860 => std_logic_vector'(x"608c0ddd"),
  1861 => std_logic_vector'(x"d17c4057"),
  1862 => std_logic_vector'(x"61104002"),
  1863 => std_logic_vector'(x"40026111"),
  1864 => std_logic_vector'(x"40c440c4"),
  1865 => std_logic_vector'(x"6110d17c"),
  1866 => std_logic_vector'(x"608c0df9"),
  1867 => std_logic_vector'(x"608c804b"),
  1868 => std_logic_vector'(x"0e85804b"),
  1869 => std_logic_vector'(x"804b608c"),
  1870 => std_logic_vector'(x"608c0e8a"),
  1871 => std_logic_vector'(x"608c8055"),
  1872 => std_logic_vector'(x"608cd1e8"),
  1873 => std_logic_vector'(x"0e8a8055"),
  1874 => std_logic_vector'(x"8055608c"),
  1875 => std_logic_vector'(x"608c0e85"),
  1876 => std_logic_vector'(x"608cd218"),
  1877 => std_logic_vector'(x"608cd22c"),
  1878 => std_logic_vector'(x"608cd240"),
  1879 => std_logic_vector'(x"608cd254"),
  1880 => std_logic_vector'(x"608cd268"),
  1881 => std_logic_vector'(x"0660d27c"),
  1882 => std_logic_vector'(x"0660d294"),
  1883 => std_logic_vector'(x"0660d2ac"),
  1884 => std_logic_vector'(x"608cd2c4"),
  1885 => std_logic_vector'(x"80018087"),
  1886 => std_logic_vector'(x"80074ea2"),
  1887 => std_logic_vector'(x"60114ea5"),
  1888 => std_logic_vector'(x"69038005"),
  1889 => std_logic_vector'(x"62038004"),
  1890 => std_logic_vector'(x"44e8d254"),
  1891 => std_logic_vector'(x"6303801f"),
  1892 => std_logic_vector'(x"6a038002"),
  1893 => std_logic_vector'(x"4ea58008"),
  1894 => std_logic_vector'(x"80066011"),
  1895 => std_logic_vector'(x"40536903"),
  1896 => std_logic_vector'(x"40026403"),
  1897 => std_logic_vector'(x"44e8d240"),
  1898 => std_logic_vector'(x"80008000"),
  1899 => std_logic_vector'(x"4153d218"),
  1900 => std_logic_vector'(x"6303803f"),
  1901 => std_logic_vector'(x"40c4d218"),
  1902 => std_logic_vector'(x"4ea58009"),
  1903 => std_logic_vector'(x"8007d218"),
  1904 => std_logic_vector'(x"40c46203"),
  1905 => std_logic_vector'(x"4ea5800a"),
  1906 => std_logic_vector'(x"8006d218"),
  1907 => std_logic_vector'(x"40c46203"),
  1908 => std_logic_vector'(x"4ea5800b"),
  1909 => std_logic_vector'(x"8005d218"),
  1910 => std_logic_vector'(x"40c46203"),
  1911 => std_logic_vector'(x"4ea5800c"),
  1912 => std_logic_vector'(x"8004d218"),
  1913 => std_logic_vector'(x"00c46203"),
  1914 => std_logic_vector'(x"fe8e608c"),
  1915 => std_logic_vector'(x"6a03800f"),
  1916 => std_logic_vector'(x"6403fcb7"),
  1917 => std_logic_vector'(x"80016600"),
  1918 => std_logic_vector'(x"4153d218"),
  1919 => std_logic_vector'(x"d2548004"),
  1920 => std_logic_vector'(x"800844e8"),
  1921 => std_logic_vector'(x"04e8d240"),
  1922 => std_logic_vector'(x"d322608c"),
  1923 => std_logic_vector'(x"d254479b"),
  1924 => std_logic_vector'(x"474f44f7"),
  1925 => std_logic_vector'(x"d32a402e"),
  1926 => std_logic_vector'(x"d240479b"),
  1927 => std_logic_vector'(x"474f44f7"),
  1928 => std_logic_vector'(x"d32e402e"),
  1929 => std_logic_vector'(x"d268479b"),
  1930 => std_logic_vector'(x"474f44f7"),
  1931 => std_logic_vector'(x"d335402e"),
  1932 => std_logic_vector'(x"d218479b"),
  1933 => std_logic_vector'(x"474b414c"),
  1934 => std_logic_vector'(x"d33c402e"),
  1935 => std_logic_vector'(x"d22c479b"),
  1936 => std_logic_vector'(x"474b414c"),
  1937 => std_logic_vector'(x"d218402e"),
  1938 => std_logic_vector'(x"d268414c"),
  1939 => std_logic_vector'(x"d25444f7"),
  1940 => std_logic_vector'(x"d24044f7"),
  1941 => std_logic_vector'(x"41c544f7"),
  1942 => std_logic_vector'(x"800146b5"),
  1943 => std_logic_vector'(x"6a03801c"),
  1944 => std_logic_vector'(x"d34241e5"),
  1945 => std_logic_vector'(x"474f479b"),
  1946 => std_logic_vector'(x"002e6103"),
  1947 => std_logic_vector'(x"d254608c"),
  1948 => std_logic_vector'(x"d24044f7"),
  1949 => std_logic_vector'(x"41aa44f7"),
  1950 => std_logic_vector'(x"4ce94eb2"),
  1951 => std_logic_vector'(x"4d304d43"),
  1952 => std_logic_vector'(x"414cd218"),
  1953 => std_logic_vector'(x"2f464d56"),
  1954 => std_logic_vector'(x"450c8084"),
  1955 => std_logic_vector'(x"44e8d268"),
  1956 => std_logic_vector'(x"80008006"),
  1957 => std_logic_vector'(x"61274448"),
  1958 => std_logic_vector'(x"44cad2c4"),
  1959 => std_logic_vector'(x"6203400b"),
  1960 => std_logic_vector'(x"d25444f7"),
  1961 => std_logic_vector'(x"800144e8"),
  1962 => std_logic_vector'(x"80008001"),
  1963 => std_logic_vector'(x"61274448"),
  1964 => std_logic_vector'(x"80806011"),
  1965 => std_logic_vector'(x"2f5e400f"),
  1966 => std_logic_vector'(x"0f7f6b1d"),
  1967 => std_logic_vector'(x"44f7d254"),
  1968 => std_logic_vector'(x"41c56111"),
  1969 => std_logic_vector'(x"47c48002"),
  1970 => std_logic_vector'(x"406441aa"),
  1971 => std_logic_vector'(x"4153d22c"),
  1972 => std_logic_vector'(x"4eb44064"),
  1973 => std_logic_vector'(x"2f6e4167"),
  1974 => std_logic_vector'(x"0f73405e"),
  1975 => std_logic_vector'(x"41674eb6"),
  1976 => std_logic_vector'(x"6b1d2f73"),
  1977 => std_logic_vector'(x"60110f7f"),
  1978 => std_logic_vector'(x"68038002"),
  1979 => std_logic_vector'(x"40022f79"),
  1980 => std_logic_vector'(x"80020f7b"),
  1981 => std_logic_vector'(x"80006203"),
  1982 => std_logic_vector'(x"44906b1d"),
  1983 => std_logic_vector'(x"43bc2f57"),
  1984 => std_logic_vector'(x"80816011"),
  1985 => std_logic_vector'(x"2f866803"),
  1986 => std_logic_vector'(x"0f8b6b1d"),
  1987 => std_logic_vector'(x"6b1d6103"),
  1988 => std_logic_vector'(x"2f8b4462"),
  1989 => std_logic_vector'(x"43bc0f4b"),
  1990 => std_logic_vector'(x"61118080"),
  1991 => std_logic_vector'(x"2f926803"),
  1992 => std_logic_vector'(x"450c8083"),
  1993 => std_logic_vector'(x"44e8d240"),
  1994 => std_logic_vector'(x"d22c6103"),
  1995 => std_logic_vector'(x"8001414c"),
  1996 => std_logic_vector'(x"6a03801c"),
  1997 => std_logic_vector'(x"44f7d268"),
  1998 => std_logic_vector'(x"d21846b5"),
  1999 => std_logic_vector'(x"608c0153"),
  2000 => std_logic_vector'(x"80108089"),
  2001 => std_logic_vector'(x"80874ea2"),
  2002 => std_logic_vector'(x"4ea28030"),
  2003 => std_logic_vector'(x"44f7d240"),
  2004 => std_logic_vector'(x"80024004"),
  2005 => std_logic_vector'(x"d2546903"),
  2006 => std_logic_vector'(x"800444f7"),
  2007 => std_logic_vector'(x"8005410a"),
  2008 => std_logic_vector'(x"64036a03"),
  2009 => std_logic_vector'(x"61108007"),
  2010 => std_logic_vector'(x"d2184ea2"),
  2011 => std_logic_vector'(x"62038004"),
  2012 => std_logic_vector'(x"800c4084"),
  2013 => std_logic_vector'(x"4ea26110"),
  2014 => std_logic_vector'(x"8005d218"),
  2015 => std_logic_vector'(x"40846203"),
  2016 => std_logic_vector'(x"6110800b"),
  2017 => std_logic_vector'(x"d2184ea2"),
  2018 => std_logic_vector'(x"62038006"),
  2019 => std_logic_vector'(x"800a4084"),
  2020 => std_logic_vector'(x"4ea26110"),
  2021 => std_logic_vector'(x"8007d218"),
  2022 => std_logic_vector'(x"40846203"),
  2023 => std_logic_vector'(x"61108009"),
  2024 => std_logic_vector'(x"d2404ea2"),
  2025 => std_logic_vector'(x"400444f7"),
  2026 => std_logic_vector'(x"6a038006"),
  2027 => std_logic_vector'(x"4084d218"),
  2028 => std_logic_vector'(x"6303803f"),
  2029 => std_logic_vector'(x"80086403"),
  2030 => std_logic_vector'(x"4ea26110"),
  2031 => std_logic_vector'(x"80008089"),
  2032 => std_logic_vector'(x"80874ea2"),
  2033 => std_logic_vector'(x"0ea28040"),
  2034 => std_logic_vector'(x"8004608c"),
  2035 => std_logic_vector'(x"80704e7a"),
  2036 => std_logic_vector'(x"d1e84ddd"),
  2037 => std_logic_vector'(x"800a44e8"),
  2038 => std_logic_vector'(x"4dc08070"),
  2039 => std_logic_vector'(x"4f374eba"),
  2040 => std_logic_vector'(x"d1e84fa0"),
  2041 => std_logic_vector'(x"807044f7"),
  2042 => std_logic_vector'(x"608c0dc0"),
  2043 => std_logic_vector'(x"608c806e"),
  2044 => std_logic_vector'(x"0e8a806e"),
  2045 => std_logic_vector'(x"806e608c"),
  2046 => std_logic_vector'(x"608c0e85"),
  2047 => std_logic_vector'(x"608cd3c0"),
  2048 => std_logic_vector'(x"608cd3d0"),
  2049 => std_logic_vector'(x"608cd3e0"),
  2050 => std_logic_vector'(x"608cd3f0"),
  2051 => std_logic_vector'(x"608cd40c"),
  2052 => std_logic_vector'(x"608cd41c"),
  2053 => std_logic_vector'(x"608cd430"),
  2054 => std_logic_vector'(x"608cd448"),
  2055 => std_logic_vector'(x"800f9954"),
  2056 => std_logic_vector'(x"fe206a03"),
  2057 => std_logic_vector'(x"608c6403"),
  2058 => std_logic_vector'(x"0660d46c"),
  2059 => std_logic_vector'(x"0660d484"),
  2060 => std_logic_vector'(x"800f8094"),
  2061 => std_logic_vector'(x"dff86a03"),
  2062 => std_logic_vector'(x"d3e06403"),
  2063 => std_logic_vector'(x"800a44e8"),
  2064 => std_logic_vector'(x"44e8d3d0"),
  2065 => std_logic_vector'(x"8001500e"),
  2066 => std_logic_vector'(x"6a038012"),
  2067 => std_logic_vector'(x"d3d041aa"),
  2068 => std_logic_vector'(x"d3e044f7"),
  2069 => std_logic_vector'(x"46b544f7"),
  2070 => std_logic_vector'(x"4153d448"),
  2071 => std_logic_vector'(x"479bd4a0"),
  2072 => std_logic_vector'(x"44f7d3e0"),
  2073 => std_logic_vector'(x"d4ad474f"),
  2074 => std_logic_vector'(x"d3d0479b"),
  2075 => std_logic_vector'(x"474f44f7"),
  2076 => std_logic_vector'(x"479bd4b5"),
  2077 => std_logic_vector'(x"414cd448"),
  2078 => std_logic_vector'(x"608c074b"),
  2079 => std_logic_vector'(x"4ffb8000"),
  2080 => std_logic_vector'(x"80066011"),
  2081 => std_logic_vector'(x"d3c06903"),
  2082 => std_logic_vector'(x"803f44e8"),
  2083 => std_logic_vector'(x"80116303"),
  2084 => std_logic_vector'(x"d3e06a03"),
  2085 => std_logic_vector'(x"800444e8"),
  2086 => std_logic_vector'(x"80094ffb"),
  2087 => std_logic_vector'(x"d3e06a03"),
  2088 => std_logic_vector'(x"640344f7"),
  2089 => std_logic_vector'(x"44e8d3e0"),
  2090 => std_logic_vector'(x"4ffb8008"),
  2091 => std_logic_vector'(x"6a038001"),
  2092 => std_logic_vector'(x"44f7d3e0"),
  2093 => std_logic_vector'(x"d3e06403"),
  2094 => std_logic_vector'(x"800c44e8"),
  2095 => std_logic_vector'(x"60114ffb"),
  2096 => std_logic_vector'(x"69038007"),
  2097 => std_logic_vector'(x"44f7d3e0"),
  2098 => std_logic_vector'(x"d3e06403"),
  2099 => std_logic_vector'(x"807f44e8"),
  2100 => std_logic_vector'(x"d3d06303"),
  2101 => std_logic_vector'(x"801444e8"),
  2102 => std_logic_vector'(x"60114ffb"),
  2103 => std_logic_vector'(x"69038006"),
  2104 => std_logic_vector'(x"6203d3f0"),
  2105 => std_logic_vector'(x"d41c4084"),
  2106 => std_logic_vector'(x"802044e8"),
  2107 => std_logic_vector'(x"80176303"),
  2108 => std_logic_vector'(x"410a8005"),
  2109 => std_logic_vector'(x"d3e06a03"),
  2110 => std_logic_vector'(x"640344f7"),
  2111 => std_logic_vector'(x"44e8d3e0"),
  2112 => std_logic_vector'(x"8001500e"),
  2113 => std_logic_vector'(x"6a038012"),
  2114 => std_logic_vector'(x"d3d041aa"),
  2115 => std_logic_vector'(x"d3e044f7"),
  2116 => std_logic_vector'(x"46b544f7"),
  2117 => std_logic_vector'(x"4153d448"),
  2118 => std_logic_vector'(x"479bd4d6"),
  2119 => std_logic_vector'(x"44f7d3e0"),
  2120 => std_logic_vector'(x"d4e3474f"),
  2121 => std_logic_vector'(x"d3d0479b"),
  2122 => std_logic_vector'(x"474f44f7"),
  2123 => std_logic_vector'(x"479bd4eb"),
  2124 => std_logic_vector'(x"414cd448"),
  2125 => std_logic_vector'(x"608c074b"),
  2126 => std_logic_vector'(x"80008004"),
  2127 => std_logic_vector'(x"61274448"),
  2128 => std_logic_vector'(x"d40c44ca"),
  2129 => std_logic_vector'(x"800244e8"),
  2130 => std_logic_vector'(x"44e8d3d0"),
  2131 => std_logic_vector'(x"80008001"),
  2132 => std_logic_vector'(x"61274448"),
  2133 => std_logic_vector'(x"d40cd3f0"),
  2134 => std_logic_vector'(x"400b44f7"),
  2135 => std_logic_vector'(x"44f76203"),
  2136 => std_logic_vector'(x"d41c6011"),
  2137 => std_logic_vector'(x"d3d044e8"),
  2138 => std_logic_vector'(x"807e44f7"),
  2139 => std_logic_vector'(x"68036111"),
  2140 => std_logic_vector'(x"610330bd"),
  2141 => std_logic_vector'(x"6b1d6103"),
  2142 => std_logic_vector'(x"467410e2"),
  2143 => std_logic_vector'(x"47c48002"),
  2144 => std_logic_vector'(x"46b58001"),
  2145 => std_logic_vector'(x"d4304064"),
  2146 => std_logic_vector'(x"40644153"),
  2147 => std_logic_vector'(x"41675014"),
  2148 => std_logic_vector'(x"405e30cb"),
  2149 => std_logic_vector'(x"501610d2"),
  2150 => std_logic_vector'(x"30d24167"),
  2151 => std_logic_vector'(x"479bd50c"),
  2152 => std_logic_vector'(x"10e26b1d"),
  2153 => std_logic_vector'(x"44f7d3d0"),
  2154 => std_logic_vector'(x"80066011"),
  2155 => std_logic_vector'(x"30da6803"),
  2156 => std_logic_vector'(x"10dc4002"),
  2157 => std_logic_vector'(x"62038002"),
  2158 => std_logic_vector'(x"44e8d3d0"),
  2159 => std_logic_vector'(x"6b1d8000"),
  2160 => std_logic_vector'(x"30a94490"),
  2161 => std_logic_vector'(x"d3d043bc"),
  2162 => std_logic_vector'(x"807f44f7"),
  2163 => std_logic_vector'(x"30ea6803"),
  2164 => std_logic_vector'(x"10ef6b1d"),
  2165 => std_logic_vector'(x"6b1d494d"),
  2166 => std_logic_vector'(x"30ef4462"),
  2167 => std_logic_vector'(x"43bc109f"),
  2168 => std_logic_vector'(x"d4306103"),
  2169 => std_logic_vector'(x"4064414c"),
  2170 => std_logic_vector'(x"479bd514"),
  2171 => std_logic_vector'(x"8001474b"),
  2172 => std_logic_vector'(x"6a038012"),
  2173 => std_logic_vector'(x"4ce98000"),
  2174 => std_logic_vector'(x"d4484d43"),
  2175 => std_logic_vector'(x"4064414c"),
  2176 => std_logic_vector'(x"479bd51a"),
  2177 => std_logic_vector'(x"4d56474b"),
  2178 => std_logic_vector'(x"800f81ff"),
  2179 => std_logic_vector'(x"ffff6a03"),
  2180 => std_logic_vector'(x"80006403"),
  2181 => std_logic_vector'(x"41674072"),
  2182 => std_logic_vector'(x"d5203112"),
  2183 => std_logic_vector'(x"474b479b"),
  2184 => std_logic_vector'(x"450c8087"),
  2185 => std_logic_vector'(x"d5354064"),
  2186 => std_logic_vector'(x"474b479b"),
  2187 => std_logic_vector'(x"d3e06103"),
  2188 => std_logic_vector'(x"608c04e8"),
  2189 => std_logic_vector'(x"44f7d3e0"),
  2190 => std_logic_vector'(x"44f7d3c0"),
  2191 => std_logic_vector'(x"6a038006"),
  2192 => std_logic_vector'(x"80fc6111"),
  2193 => std_logic_vector'(x"6a03800f"),
  2194 => std_logic_vector'(x"64038000"),
  2195 => std_logic_vector'(x"80116303"),
  2196 => std_logic_vector'(x"64036903"),
  2197 => std_logic_vector'(x"61108003"),
  2198 => std_logic_vector'(x"60114ff8"),
  2199 => std_logic_vector'(x"69038009"),
  2200 => std_logic_vector'(x"630380ff"),
  2201 => std_logic_vector'(x"61108007"),
  2202 => std_logic_vector'(x"60114ff8"),
  2203 => std_logic_vector'(x"69038001"),
  2204 => std_logic_vector'(x"630380ff"),
  2205 => std_logic_vector'(x"6110800b"),
  2206 => std_logic_vector'(x"60114ff8"),
  2207 => std_logic_vector'(x"63038001"),
  2208 => std_logic_vector'(x"6a038007"),
  2209 => std_logic_vector'(x"44f7d3d0"),
  2210 => std_logic_vector'(x"6303807f"),
  2211 => std_logic_vector'(x"800f6403"),
  2212 => std_logic_vector'(x"4ff86110"),
  2213 => std_logic_vector'(x"4ffb8014"),
  2214 => std_logic_vector'(x"6303801f"),
  2215 => std_logic_vector'(x"44f7d40c"),
  2216 => std_logic_vector'(x"6a038006"),
  2217 => std_logic_vector'(x"61106403"),
  2218 => std_logic_vector'(x"800f8018"),
  2219 => std_logic_vector'(x"b5006a03"),
  2220 => std_logic_vector'(x"63036403"),
  2221 => std_logic_vector'(x"80058017"),
  2222 => std_logic_vector'(x"6903410a"),
  2223 => std_logic_vector'(x"80176403"),
  2224 => std_logic_vector'(x"4ff86110"),
  2225 => std_logic_vector'(x"4ffb8012"),
  2226 => std_logic_vector'(x"80e76011"),
  2227 => std_logic_vector'(x"80126303"),
  2228 => std_logic_vector'(x"4ff86110"),
  2229 => std_logic_vector'(x"64038018"),
  2230 => std_logic_vector'(x"61108012"),
  2231 => std_logic_vector'(x"608c0ff8"),
  2232 => std_logic_vector'(x"509c503e"),
  2233 => std_logic_vector'(x"608c111a"),
  2234 => std_logic_vector'(x"80006111"),
  2235 => std_logic_vector'(x"68036600"),
  2236 => std_logic_vector'(x"47c48002"),
  2237 => std_logic_vector'(x"400f800f"),
  2238 => std_logic_vector'(x"31826403"),
  2239 => std_logic_vector'(x"479bd574"),
  2240 => std_logic_vector'(x"450c8083"),
  2241 => std_logic_vector'(x"80006011"),
  2242 => std_logic_vector'(x"61116803"),
  2243 => std_logic_vector'(x"400f800f"),
  2244 => std_logic_vector'(x"318e6403"),
  2245 => std_logic_vector'(x"479bd594"),
  2246 => std_logic_vector'(x"450c8083"),
  2247 => std_logic_vector'(x"4e7a8004"),
  2248 => std_logic_vector'(x"4ddd8070"),
  2249 => std_logic_vector'(x"44e8d1e8"),
  2250 => std_logic_vector'(x"8070800c"),
  2251 => std_logic_vector'(x"61114dc0"),
  2252 => std_logic_vector'(x"66008000"),
  2253 => std_logic_vector'(x"31a26703"),
  2254 => std_logic_vector'(x"62038020"),
  2255 => std_logic_vector'(x"4e9b8000"),
  2256 => std_logic_vector'(x"11c76103"),
  2257 => std_logic_vector'(x"80016011"),
  2258 => std_logic_vector'(x"31ab6303"),
  2259 => std_logic_vector'(x"80046110"),
  2260 => std_logic_vector'(x"800f6a03"),
  2261 => std_logic_vector'(x"611011ad"),
  2262 => std_logic_vector'(x"405380f0"),
  2263 => std_logic_vector'(x"61276011"),
  2264 => std_logic_vector'(x"69038001"),
  2265 => std_logic_vector'(x"62038090"),
  2266 => std_logic_vector'(x"6b116127"),
  2267 => std_logic_vector'(x"63034e98"),
  2268 => std_logic_vector'(x"6b1d6403"),
  2269 => std_logic_vector'(x"4e9b6110"),
  2270 => std_logic_vector'(x"80008081"),
  2271 => std_logic_vector'(x"80804e9b"),
  2272 => std_logic_vector'(x"4e9b8001"),
  2273 => std_logic_vector'(x"80206b1d"),
  2274 => std_logic_vector'(x"80306203"),
  2275 => std_logic_vector'(x"d1e84e9b"),
  2276 => std_logic_vector'(x"807044f7"),
  2277 => std_logic_vector'(x"608c0dc0"),
  2278 => std_logic_vector'(x"608cd5c0"),
  2279 => std_logic_vector'(x"608c8058"),
  2280 => std_logic_vector'(x"608c800c"),
  2281 => std_logic_vector'(x"4e7a8004"),
  2282 => std_logic_vector'(x"8070800c"),
  2283 => std_logic_vector'(x"80984dc0"),
  2284 => std_logic_vector'(x"4dc08058"),
  2285 => std_logic_vector'(x"8008d5c0"),
  2286 => std_logic_vector'(x"0e268058"),
  2287 => std_logic_vector'(x"8000608c"),
  2288 => std_logic_vector'(x"61274448"),
  2289 => std_logic_vector'(x"44ca6011"),
  2290 => std_logic_vector'(x"40846203"),
  2291 => std_logic_vector'(x"6b1d474f"),
  2292 => std_logic_vector'(x"31eb4462"),
  2293 => std_logic_vector'(x"43bc11e1"),
  2294 => std_logic_vector'(x"608c6103"),
  2295 => std_logic_vector'(x"4e7a8004"),
  2296 => std_logic_vector'(x"80704d97"),
  2297 => std_logic_vector'(x"074f4ddd"),
  2298 => std_logic_vector'(x"0000608c"),
  2299 => std_logic_vector'(x"00000000"),
  2300 => std_logic_vector'(x"00000000"),
  2301 => std_logic_vector'(x"00000000"),
  2302 => std_logic_vector'(x"00000000"),
  2303 => std_logic_vector'(x"00000000"),
  2304 => std_logic_vector'(x"00000000"),
  2305 => std_logic_vector'(x"00000000"),
  2306 => std_logic_vector'(x"00000000"),
  2307 => std_logic_vector'(x"00000000"),
  2308 => std_logic_vector'(x"00000000"),
  2309 => std_logic_vector'(x"00000000"),
  2310 => std_logic_vector'(x"00000000"),
  2311 => std_logic_vector'(x"00000000"),
  2312 => std_logic_vector'(x"00000000"),
  2313 => std_logic_vector'(x"00000000"),
  2314 => std_logic_vector'(x"00000000"),
  2315 => std_logic_vector'(x"00000000"),
  2316 => std_logic_vector'(x"00000000"),
  2317 => std_logic_vector'(x"00000000"),
  2318 => std_logic_vector'(x"00000000"),
  2319 => std_logic_vector'(x"00000000"),
  2320 => std_logic_vector'(x"00000000"),
  2321 => std_logic_vector'(x"00000000"),
  2322 => std_logic_vector'(x"00000000"),
  2323 => std_logic_vector'(x"00000000"),
  2324 => std_logic_vector'(x"00000000"),
  2325 => std_logic_vector'(x"00000000"),
  2326 => std_logic_vector'(x"00000000"),
  2327 => std_logic_vector'(x"00000000"),
  2328 => std_logic_vector'(x"00000000"),
  2329 => std_logic_vector'(x"00000000"),
  2330 => std_logic_vector'(x"00000000"),
  2331 => std_logic_vector'(x"00000000"),
  2332 => std_logic_vector'(x"00000000"),
  2333 => std_logic_vector'(x"00000000"),
  2334 => std_logic_vector'(x"00000000"),
  2335 => std_logic_vector'(x"00000000"),
  2336 => std_logic_vector'(x"00000000"),
  2337 => std_logic_vector'(x"00000000"),
  2338 => std_logic_vector'(x"00000000"),
  2339 => std_logic_vector'(x"00000000"),
  2340 => std_logic_vector'(x"00000000"),
  2341 => std_logic_vector'(x"00000000"),
  2342 => std_logic_vector'(x"00000000"),
  2343 => std_logic_vector'(x"00000000"),
  2344 => std_logic_vector'(x"00000000"),
  2345 => std_logic_vector'(x"00000000"),
  2346 => std_logic_vector'(x"00000000"),
  2347 => std_logic_vector'(x"00000000"),
  2348 => std_logic_vector'(x"00000000"),
  2349 => std_logic_vector'(x"00000000"),
  2350 => std_logic_vector'(x"00000000"),
  2351 => std_logic_vector'(x"00000000"),
  2352 => std_logic_vector'(x"00000000"),
  2353 => std_logic_vector'(x"00000000"),
  2354 => std_logic_vector'(x"00000000"),
  2355 => std_logic_vector'(x"00000000"),
  2356 => std_logic_vector'(x"00000000"),
  2357 => std_logic_vector'(x"00000000"),
  2358 => std_logic_vector'(x"00000000"),
  2359 => std_logic_vector'(x"00000000"),
  2360 => std_logic_vector'(x"00000000"),
  2361 => std_logic_vector'(x"00000000"),
  2362 => std_logic_vector'(x"00000000"),
  2363 => std_logic_vector'(x"00000000"),
  2364 => std_logic_vector'(x"00000000"),
  2365 => std_logic_vector'(x"00000000"),
  2366 => std_logic_vector'(x"00000000"),
  2367 => std_logic_vector'(x"00000000"),
  2368 => std_logic_vector'(x"00000000"),
  2369 => std_logic_vector'(x"00000000"),
  2370 => std_logic_vector'(x"00000000"),
  2371 => std_logic_vector'(x"00000000"),
  2372 => std_logic_vector'(x"00000000"),
  2373 => std_logic_vector'(x"00000000"),
  2374 => std_logic_vector'(x"00000000"),
  2375 => std_logic_vector'(x"00000000"),
  2376 => std_logic_vector'(x"00000000"),
  2377 => std_logic_vector'(x"00000000"),
  2378 => std_logic_vector'(x"00000000"),
  2379 => std_logic_vector'(x"00000000"),
  2380 => std_logic_vector'(x"00000000"),
  2381 => std_logic_vector'(x"00000000"),
  2382 => std_logic_vector'(x"00000000"),
  2383 => std_logic_vector'(x"00000000"),
  2384 => std_logic_vector'(x"00000000"),
  2385 => std_logic_vector'(x"00000000"),
  2386 => std_logic_vector'(x"00000000"),
  2387 => std_logic_vector'(x"00000000"),
  2388 => std_logic_vector'(x"00000000"),
  2389 => std_logic_vector'(x"00000000"),
  2390 => std_logic_vector'(x"00000000"),
  2391 => std_logic_vector'(x"00000000"),
  2392 => std_logic_vector'(x"00000000"),
  2393 => std_logic_vector'(x"00000000"),
  2394 => std_logic_vector'(x"00000000"),
  2395 => std_logic_vector'(x"00000000"),
  2396 => std_logic_vector'(x"00000000"),
  2397 => std_logic_vector'(x"00000000"),
  2398 => std_logic_vector'(x"00000000"),
  2399 => std_logic_vector'(x"00000000"),
  2400 => std_logic_vector'(x"00000000"),
  2401 => std_logic_vector'(x"00000000"),
  2402 => std_logic_vector'(x"00000000"),
  2403 => std_logic_vector'(x"00000000"),
  2404 => std_logic_vector'(x"00000000"),
  2405 => std_logic_vector'(x"00000000"),
  2406 => std_logic_vector'(x"00000000"),
  2407 => std_logic_vector'(x"00000000"),
  2408 => std_logic_vector'(x"00000000"),
  2409 => std_logic_vector'(x"00000000"),
  2410 => std_logic_vector'(x"00000000"),
  2411 => std_logic_vector'(x"00000000"),
  2412 => std_logic_vector'(x"00000000"),
  2413 => std_logic_vector'(x"00000000"),
  2414 => std_logic_vector'(x"00000000"),
  2415 => std_logic_vector'(x"00000000"),
  2416 => std_logic_vector'(x"00000000"),
  2417 => std_logic_vector'(x"00000000"),
  2418 => std_logic_vector'(x"00000000"),
  2419 => std_logic_vector'(x"00000000"),
  2420 => std_logic_vector'(x"00000000"),
  2421 => std_logic_vector'(x"00000000"),
  2422 => std_logic_vector'(x"00000000"),
  2423 => std_logic_vector'(x"00000000"),
  2424 => std_logic_vector'(x"00000000"),
  2425 => std_logic_vector'(x"00000000"),
  2426 => std_logic_vector'(x"00000000"),
  2427 => std_logic_vector'(x"00000000"),
  2428 => std_logic_vector'(x"00000000"),
  2429 => std_logic_vector'(x"00000000"),
  2430 => std_logic_vector'(x"00000000"),
  2431 => std_logic_vector'(x"00000000"),
  2432 => std_logic_vector'(x"00000000"),
  2433 => std_logic_vector'(x"00000000"),
  2434 => std_logic_vector'(x"00000000"),
  2435 => std_logic_vector'(x"00000000"),
  2436 => std_logic_vector'(x"00000000"),
  2437 => std_logic_vector'(x"00000000"),
  2438 => std_logic_vector'(x"00000000"),
  2439 => std_logic_vector'(x"00000000"),
  2440 => std_logic_vector'(x"00000000"),
  2441 => std_logic_vector'(x"00000000"),
  2442 => std_logic_vector'(x"00000000"),
  2443 => std_logic_vector'(x"00000000"),
  2444 => std_logic_vector'(x"00000000"),
  2445 => std_logic_vector'(x"00000000"),
  2446 => std_logic_vector'(x"00000000"),
  2447 => std_logic_vector'(x"00000000"),
  2448 => std_logic_vector'(x"00000000"),
  2449 => std_logic_vector'(x"00000000"),
  2450 => std_logic_vector'(x"00000000"),
  2451 => std_logic_vector'(x"00000000"),
  2452 => std_logic_vector'(x"00000000"),
  2453 => std_logic_vector'(x"00000000"),
  2454 => std_logic_vector'(x"00000000"),
  2455 => std_logic_vector'(x"00000000"),
  2456 => std_logic_vector'(x"00000000"),
  2457 => std_logic_vector'(x"00000000"),
  2458 => std_logic_vector'(x"00000000"),
  2459 => std_logic_vector'(x"00000000"),
  2460 => std_logic_vector'(x"00000000"),
  2461 => std_logic_vector'(x"00000000"),
  2462 => std_logic_vector'(x"00000000"),
  2463 => std_logic_vector'(x"00000000"),
  2464 => std_logic_vector'(x"00000000"),
  2465 => std_logic_vector'(x"00000000"),
  2466 => std_logic_vector'(x"00000000"),
  2467 => std_logic_vector'(x"00000000"),
  2468 => std_logic_vector'(x"00000000"),
  2469 => std_logic_vector'(x"00000000"),
  2470 => std_logic_vector'(x"00000000"),
  2471 => std_logic_vector'(x"00000000"),
  2472 => std_logic_vector'(x"00000000"),
  2473 => std_logic_vector'(x"00000000"),
  2474 => std_logic_vector'(x"00000000"),
  2475 => std_logic_vector'(x"00000000"),
  2476 => std_logic_vector'(x"00000000"),
  2477 => std_logic_vector'(x"00000000"),
  2478 => std_logic_vector'(x"00000000"),
  2479 => std_logic_vector'(x"00000000"),
  2480 => std_logic_vector'(x"00000000"),
  2481 => std_logic_vector'(x"00000000"),
  2482 => std_logic_vector'(x"00000000"),
  2483 => std_logic_vector'(x"00000000"),
  2484 => std_logic_vector'(x"00000000"),
  2485 => std_logic_vector'(x"00000000"),
  2486 => std_logic_vector'(x"00000000"),
  2487 => std_logic_vector'(x"00000000"),
  2488 => std_logic_vector'(x"00000000"),
  2489 => std_logic_vector'(x"00000000"),
  2490 => std_logic_vector'(x"00000000"),
  2491 => std_logic_vector'(x"00000000"),
  2492 => std_logic_vector'(x"00000000"),
  2493 => std_logic_vector'(x"00000000"),
  2494 => std_logic_vector'(x"00000000"),
  2495 => std_logic_vector'(x"00000000"),
  2496 => std_logic_vector'(x"00000000"),
  2497 => std_logic_vector'(x"00000000"),
  2498 => std_logic_vector'(x"00000000"),
  2499 => std_logic_vector'(x"00000000"),
  2500 => std_logic_vector'(x"00000000"),
  2501 => std_logic_vector'(x"00000000"),
  2502 => std_logic_vector'(x"00000000"),
  2503 => std_logic_vector'(x"00000000"),
  2504 => std_logic_vector'(x"00000000"),
  2505 => std_logic_vector'(x"00000000"),
  2506 => std_logic_vector'(x"00000000"),
  2507 => std_logic_vector'(x"00000000"),
  2508 => std_logic_vector'(x"00000000"),
  2509 => std_logic_vector'(x"00000000"),
  2510 => std_logic_vector'(x"00000000"),
  2511 => std_logic_vector'(x"00000000"),
  2512 => std_logic_vector'(x"00000000"),
  2513 => std_logic_vector'(x"00000000"),
  2514 => std_logic_vector'(x"00000000"),
  2515 => std_logic_vector'(x"00000000"),
  2516 => std_logic_vector'(x"00000000"),
  2517 => std_logic_vector'(x"00000000"),
  2518 => std_logic_vector'(x"00000000"),
  2519 => std_logic_vector'(x"00000000"),
  2520 => std_logic_vector'(x"00000000"),
  2521 => std_logic_vector'(x"00000000"),
  2522 => std_logic_vector'(x"00000000"),
  2523 => std_logic_vector'(x"00000000"),
  2524 => std_logic_vector'(x"00000000"),
  2525 => std_logic_vector'(x"00000000"),
  2526 => std_logic_vector'(x"00000000"),
  2527 => std_logic_vector'(x"00000000"),
  2528 => std_logic_vector'(x"00000000"),
  2529 => std_logic_vector'(x"00000000"),
  2530 => std_logic_vector'(x"00000000"),
  2531 => std_logic_vector'(x"00000000"),
  2532 => std_logic_vector'(x"00000000"),
  2533 => std_logic_vector'(x"00000000"),
  2534 => std_logic_vector'(x"00000000"),
  2535 => std_logic_vector'(x"00000000"),
  2536 => std_logic_vector'(x"00000000"),
  2537 => std_logic_vector'(x"00000000"),
  2538 => std_logic_vector'(x"00000000"),
  2539 => std_logic_vector'(x"00000000"),
  2540 => std_logic_vector'(x"00000000"),
  2541 => std_logic_vector'(x"00000000"),
  2542 => std_logic_vector'(x"00000000"),
  2543 => std_logic_vector'(x"00000000"),
  2544 => std_logic_vector'(x"00000000"),
  2545 => std_logic_vector'(x"00000000"),
  2546 => std_logic_vector'(x"00000000"),
  2547 => std_logic_vector'(x"00000000"),
  2548 => std_logic_vector'(x"00000000"),
  2549 => std_logic_vector'(x"00000000"),
  2550 => std_logic_vector'(x"00000000"),
  2551 => std_logic_vector'(x"00000000"),
  2552 => std_logic_vector'(x"00000000"),
  2553 => std_logic_vector'(x"00000000"),
  2554 => std_logic_vector'(x"00000000"),
  2555 => std_logic_vector'(x"00000000"),
  2556 => std_logic_vector'(x"00000000"),
  2557 => std_logic_vector'(x"00000000"),
  2558 => std_logic_vector'(x"00000000"),
  2559 => std_logic_vector'(x"00000000"),
  2560 => std_logic_vector'(x"00000000"),
  2561 => std_logic_vector'(x"00000000"),
  2562 => std_logic_vector'(x"00000000"),
  2563 => std_logic_vector'(x"00000000"),
  2564 => std_logic_vector'(x"00000000"),
  2565 => std_logic_vector'(x"00000000"),
  2566 => std_logic_vector'(x"00000000"),
  2567 => std_logic_vector'(x"00000000"),
  2568 => std_logic_vector'(x"00000000"),
  2569 => std_logic_vector'(x"00000000"),
  2570 => std_logic_vector'(x"00000000"),
  2571 => std_logic_vector'(x"00000000"),
  2572 => std_logic_vector'(x"00000000"),
  2573 => std_logic_vector'(x"00000000"),
  2574 => std_logic_vector'(x"00000000"),
  2575 => std_logic_vector'(x"00000000"),
  2576 => std_logic_vector'(x"00000000"),
  2577 => std_logic_vector'(x"00000000"),
  2578 => std_logic_vector'(x"00000000"),
  2579 => std_logic_vector'(x"00000000"),
  2580 => std_logic_vector'(x"00000000"),
  2581 => std_logic_vector'(x"00000000"),
  2582 => std_logic_vector'(x"00000000"),
  2583 => std_logic_vector'(x"00000000"),
  2584 => std_logic_vector'(x"00000000"),
  2585 => std_logic_vector'(x"00000000"),
  2586 => std_logic_vector'(x"00000000"),
  2587 => std_logic_vector'(x"00000000"),
  2588 => std_logic_vector'(x"00000000"),
  2589 => std_logic_vector'(x"00000000"),
  2590 => std_logic_vector'(x"00000000"),
  2591 => std_logic_vector'(x"00000000"),
  2592 => std_logic_vector'(x"00000000"),
  2593 => std_logic_vector'(x"00000000"),
  2594 => std_logic_vector'(x"00000000"),
  2595 => std_logic_vector'(x"00000000"),
  2596 => std_logic_vector'(x"00000000"),
  2597 => std_logic_vector'(x"00000000"),
  2598 => std_logic_vector'(x"00000000"),
  2599 => std_logic_vector'(x"00000000"),
  2600 => std_logic_vector'(x"00000000"),
  2601 => std_logic_vector'(x"00000000"),
  2602 => std_logic_vector'(x"00000000"),
  2603 => std_logic_vector'(x"00000000"),
  2604 => std_logic_vector'(x"00000000"),
  2605 => std_logic_vector'(x"00000000"),
  2606 => std_logic_vector'(x"00000000"),
  2607 => std_logic_vector'(x"00000000"),
  2608 => std_logic_vector'(x"00000000"),
  2609 => std_logic_vector'(x"00000000"),
  2610 => std_logic_vector'(x"00000000"),
  2611 => std_logic_vector'(x"00000000"),
  2612 => std_logic_vector'(x"00000000"),
  2613 => std_logic_vector'(x"00000000"),
  2614 => std_logic_vector'(x"00000000"),
  2615 => std_logic_vector'(x"00000000"),
  2616 => std_logic_vector'(x"00000000"),
  2617 => std_logic_vector'(x"00000000"),
  2618 => std_logic_vector'(x"00000000"),
  2619 => std_logic_vector'(x"00000000"),
  2620 => std_logic_vector'(x"00000000"),
  2621 => std_logic_vector'(x"00000000"),
  2622 => std_logic_vector'(x"00000000"),
  2623 => std_logic_vector'(x"00000000"),
  2624 => std_logic_vector'(x"00000000"),
  2625 => std_logic_vector'(x"00000000"),
  2626 => std_logic_vector'(x"00000000"),
  2627 => std_logic_vector'(x"00000000"),
  2628 => std_logic_vector'(x"00000000"),
  2629 => std_logic_vector'(x"00000000"),
  2630 => std_logic_vector'(x"00000000"),
  2631 => std_logic_vector'(x"00000000"),
  2632 => std_logic_vector'(x"00000000"),
  2633 => std_logic_vector'(x"00000000"),
  2634 => std_logic_vector'(x"00000000"),
  2635 => std_logic_vector'(x"00000000"),
  2636 => std_logic_vector'(x"00000000"),
  2637 => std_logic_vector'(x"00000000"),
  2638 => std_logic_vector'(x"00000000"),
  2639 => std_logic_vector'(x"00000000"),
  2640 => std_logic_vector'(x"00000000"),
  2641 => std_logic_vector'(x"00000000"),
  2642 => std_logic_vector'(x"00000000"),
  2643 => std_logic_vector'(x"00000000"),
  2644 => std_logic_vector'(x"00000000"),
  2645 => std_logic_vector'(x"00000000"),
  2646 => std_logic_vector'(x"00000000"),
  2647 => std_logic_vector'(x"00000000"),
  2648 => std_logic_vector'(x"00000000"),
  2649 => std_logic_vector'(x"00000000"),
  2650 => std_logic_vector'(x"00000000"),
  2651 => std_logic_vector'(x"00000000"),
  2652 => std_logic_vector'(x"00000000"),
  2653 => std_logic_vector'(x"00000000"),
  2654 => std_logic_vector'(x"00000000"),
  2655 => std_logic_vector'(x"00000000"),
  2656 => std_logic_vector'(x"00000000"),
  2657 => std_logic_vector'(x"00000000"),
  2658 => std_logic_vector'(x"00000000"),
  2659 => std_logic_vector'(x"00000000"),
  2660 => std_logic_vector'(x"00000000"),
  2661 => std_logic_vector'(x"00000000"),
  2662 => std_logic_vector'(x"00000000"),
  2663 => std_logic_vector'(x"00000000"),
  2664 => std_logic_vector'(x"00000000"),
  2665 => std_logic_vector'(x"00000000"),
  2666 => std_logic_vector'(x"00000000"),
  2667 => std_logic_vector'(x"00000000"),
  2668 => std_logic_vector'(x"00000000"),
  2669 => std_logic_vector'(x"00000000"),
  2670 => std_logic_vector'(x"00000000"),
  2671 => std_logic_vector'(x"00000000"),
  2672 => std_logic_vector'(x"00000000"),
  2673 => std_logic_vector'(x"00000000"),
  2674 => std_logic_vector'(x"00000000"),
  2675 => std_logic_vector'(x"00000000"),
  2676 => std_logic_vector'(x"00000000"),
  2677 => std_logic_vector'(x"00000000"),
  2678 => std_logic_vector'(x"00000000"),
  2679 => std_logic_vector'(x"00000000"),
  2680 => std_logic_vector'(x"00000000"),
  2681 => std_logic_vector'(x"00000000"),
  2682 => std_logic_vector'(x"00000000"),
  2683 => std_logic_vector'(x"00000000"),
  2684 => std_logic_vector'(x"00000000"),
  2685 => std_logic_vector'(x"00000000"),
  2686 => std_logic_vector'(x"00000000"),
  2687 => std_logic_vector'(x"00000000"),
  2688 => std_logic_vector'(x"00000000"),
  2689 => std_logic_vector'(x"00000000"),
  2690 => std_logic_vector'(x"00000000"),
  2691 => std_logic_vector'(x"00000000"),
  2692 => std_logic_vector'(x"00000000"),
  2693 => std_logic_vector'(x"00000000"),
  2694 => std_logic_vector'(x"00000000"),
  2695 => std_logic_vector'(x"00000000"),
  2696 => std_logic_vector'(x"00000000"),
  2697 => std_logic_vector'(x"00000000"),
  2698 => std_logic_vector'(x"00000000"),
  2699 => std_logic_vector'(x"00000000"),
  2700 => std_logic_vector'(x"00000000"),
  2701 => std_logic_vector'(x"00000000"),
  2702 => std_logic_vector'(x"00000000"),
  2703 => std_logic_vector'(x"00000000"),
  2704 => std_logic_vector'(x"00000000"),
  2705 => std_logic_vector'(x"00000000"),
  2706 => std_logic_vector'(x"00000000"),
  2707 => std_logic_vector'(x"00000000"),
  2708 => std_logic_vector'(x"00000000"),
  2709 => std_logic_vector'(x"00000000"),
  2710 => std_logic_vector'(x"00000000"),
  2711 => std_logic_vector'(x"00000000"),
  2712 => std_logic_vector'(x"00000000"),
  2713 => std_logic_vector'(x"00000000"),
  2714 => std_logic_vector'(x"00000000"),
  2715 => std_logic_vector'(x"00000000"),
  2716 => std_logic_vector'(x"00000000"),
  2717 => std_logic_vector'(x"00000000"),
  2718 => std_logic_vector'(x"00000000"),
  2719 => std_logic_vector'(x"00000000"),
  2720 => std_logic_vector'(x"00000000"),
  2721 => std_logic_vector'(x"00000000"),
  2722 => std_logic_vector'(x"00000000"),
  2723 => std_logic_vector'(x"00000000"),
  2724 => std_logic_vector'(x"00000000"),
  2725 => std_logic_vector'(x"00000000"),
  2726 => std_logic_vector'(x"00000000"),
  2727 => std_logic_vector'(x"00000000"),
  2728 => std_logic_vector'(x"00000000"),
  2729 => std_logic_vector'(x"00000000"),
  2730 => std_logic_vector'(x"00000000"),
  2731 => std_logic_vector'(x"00000000"),
  2732 => std_logic_vector'(x"00000000"),
  2733 => std_logic_vector'(x"00000000"),
  2734 => std_logic_vector'(x"00000000"),
  2735 => std_logic_vector'(x"00000000"),
  2736 => std_logic_vector'(x"00000000"),
  2737 => std_logic_vector'(x"00000000"),
  2738 => std_logic_vector'(x"00000000"),
  2739 => std_logic_vector'(x"00000000"),
  2740 => std_logic_vector'(x"00000000"),
  2741 => std_logic_vector'(x"00000000"),
  2742 => std_logic_vector'(x"00000000"),
  2743 => std_logic_vector'(x"00000000"),
  2744 => std_logic_vector'(x"00000000"),
  2745 => std_logic_vector'(x"00000000"),
  2746 => std_logic_vector'(x"00000000"),
  2747 => std_logic_vector'(x"00000000"),
  2748 => std_logic_vector'(x"00000000"),
  2749 => std_logic_vector'(x"00000000"),
  2750 => std_logic_vector'(x"00000000"),
  2751 => std_logic_vector'(x"00000000"),
  2752 => std_logic_vector'(x"00000000"),
  2753 => std_logic_vector'(x"00000000"),
  2754 => std_logic_vector'(x"00000000"),
  2755 => std_logic_vector'(x"00000000"),
  2756 => std_logic_vector'(x"00000000"),
  2757 => std_logic_vector'(x"00000000"),
  2758 => std_logic_vector'(x"00000000"),
  2759 => std_logic_vector'(x"00000000"),
  2760 => std_logic_vector'(x"00000000"),
  2761 => std_logic_vector'(x"00000000"),
  2762 => std_logic_vector'(x"00000000"),
  2763 => std_logic_vector'(x"00000000"),
  2764 => std_logic_vector'(x"00000000"),
  2765 => std_logic_vector'(x"00000000"),
  2766 => std_logic_vector'(x"00000000"),
  2767 => std_logic_vector'(x"00000000"),
  2768 => std_logic_vector'(x"00000000"),
  2769 => std_logic_vector'(x"00000000"),
  2770 => std_logic_vector'(x"00000000"),
  2771 => std_logic_vector'(x"00000000"),
  2772 => std_logic_vector'(x"00000000"),
  2773 => std_logic_vector'(x"00000000"),
  2774 => std_logic_vector'(x"00000000"),
  2775 => std_logic_vector'(x"00000000"),
  2776 => std_logic_vector'(x"00000000"),
  2777 => std_logic_vector'(x"00000000"),
  2778 => std_logic_vector'(x"00000000"),
  2779 => std_logic_vector'(x"00000000"),
  2780 => std_logic_vector'(x"00000000"),
  2781 => std_logic_vector'(x"00000000"),
  2782 => std_logic_vector'(x"00000000"),
  2783 => std_logic_vector'(x"00000000"),
  2784 => std_logic_vector'(x"00000000"),
  2785 => std_logic_vector'(x"00000000"),
  2786 => std_logic_vector'(x"00000000"),
  2787 => std_logic_vector'(x"00000000"),
  2788 => std_logic_vector'(x"00000000"),
  2789 => std_logic_vector'(x"00000000"),
  2790 => std_logic_vector'(x"00000000"),
  2791 => std_logic_vector'(x"00000000"),
  2792 => std_logic_vector'(x"00000000"),
  2793 => std_logic_vector'(x"00000000"),
  2794 => std_logic_vector'(x"00000000"),
  2795 => std_logic_vector'(x"00000000"),
  2796 => std_logic_vector'(x"00000000"),
  2797 => std_logic_vector'(x"00000000"),
  2798 => std_logic_vector'(x"00000000"),
  2799 => std_logic_vector'(x"00000000"),
  2800 => std_logic_vector'(x"00000000"),
  2801 => std_logic_vector'(x"00000000"),
  2802 => std_logic_vector'(x"00000000"),
  2803 => std_logic_vector'(x"00000000"),
  2804 => std_logic_vector'(x"00000000"),
  2805 => std_logic_vector'(x"00000000"),
  2806 => std_logic_vector'(x"00000000"),
  2807 => std_logic_vector'(x"00000000"),
  2808 => std_logic_vector'(x"00000000"),
  2809 => std_logic_vector'(x"00000000"),
  2810 => std_logic_vector'(x"00000000"),
  2811 => std_logic_vector'(x"00000000"),
  2812 => std_logic_vector'(x"00000000"),
  2813 => std_logic_vector'(x"00000000"),
  2814 => std_logic_vector'(x"00000000"),
  2815 => std_logic_vector'(x"00000000"),
  2816 => std_logic_vector'(x"00000000"),
  2817 => std_logic_vector'(x"00000000"),
  2818 => std_logic_vector'(x"00000000"),
  2819 => std_logic_vector'(x"00000000"),
  2820 => std_logic_vector'(x"00000000"),
  2821 => std_logic_vector'(x"00000000"),
  2822 => std_logic_vector'(x"00000000"),
  2823 => std_logic_vector'(x"00000000"),
  2824 => std_logic_vector'(x"00000000"),
  2825 => std_logic_vector'(x"00000000"),
  2826 => std_logic_vector'(x"00000000"),
  2827 => std_logic_vector'(x"00000000"),
  2828 => std_logic_vector'(x"00000000"),
  2829 => std_logic_vector'(x"00000000"),
  2830 => std_logic_vector'(x"00000000"),
  2831 => std_logic_vector'(x"00000000"),
  2832 => std_logic_vector'(x"00000000"),
  2833 => std_logic_vector'(x"00000000"),
  2834 => std_logic_vector'(x"00000000"),
  2835 => std_logic_vector'(x"00000000"),
  2836 => std_logic_vector'(x"00000000"),
  2837 => std_logic_vector'(x"00000000"),
  2838 => std_logic_vector'(x"00000000"),
  2839 => std_logic_vector'(x"00000000"),
  2840 => std_logic_vector'(x"00000000"),
  2841 => std_logic_vector'(x"00000000"),
  2842 => std_logic_vector'(x"00000000"),
  2843 => std_logic_vector'(x"00000000"),
  2844 => std_logic_vector'(x"00000000"),
  2845 => std_logic_vector'(x"00000000"),
  2846 => std_logic_vector'(x"00000000"),
  2847 => std_logic_vector'(x"00000000"),
  2848 => std_logic_vector'(x"00000000"),
  2849 => std_logic_vector'(x"00000000"),
  2850 => std_logic_vector'(x"00000000"),
  2851 => std_logic_vector'(x"00000000"),
  2852 => std_logic_vector'(x"00000000"),
  2853 => std_logic_vector'(x"00000000"),
  2854 => std_logic_vector'(x"00000000"),
  2855 => std_logic_vector'(x"00000000"),
  2856 => std_logic_vector'(x"00000000"),
  2857 => std_logic_vector'(x"00000000"),
  2858 => std_logic_vector'(x"00000000"),
  2859 => std_logic_vector'(x"00000000"),
  2860 => std_logic_vector'(x"00000000"),
  2861 => std_logic_vector'(x"00000000"),
  2862 => std_logic_vector'(x"00000000"),
  2863 => std_logic_vector'(x"00000000"),
  2864 => std_logic_vector'(x"00000000"),
  2865 => std_logic_vector'(x"00000000"),
  2866 => std_logic_vector'(x"00000000"),
  2867 => std_logic_vector'(x"00000000"),
  2868 => std_logic_vector'(x"00000000"),
  2869 => std_logic_vector'(x"00000000"),
  2870 => std_logic_vector'(x"00000000"),
  2871 => std_logic_vector'(x"00000000"),
  2872 => std_logic_vector'(x"00000000"),
  2873 => std_logic_vector'(x"00000000"),
  2874 => std_logic_vector'(x"00000000"),
  2875 => std_logic_vector'(x"00000000"),
  2876 => std_logic_vector'(x"00000000"),
  2877 => std_logic_vector'(x"00000000"),
  2878 => std_logic_vector'(x"00000000"),
  2879 => std_logic_vector'(x"00000000"),
  2880 => std_logic_vector'(x"00000000"),
  2881 => std_logic_vector'(x"00000000"),
  2882 => std_logic_vector'(x"00000000"),
  2883 => std_logic_vector'(x"00000000"),
  2884 => std_logic_vector'(x"00000000"),
  2885 => std_logic_vector'(x"00000000"),
  2886 => std_logic_vector'(x"00000000"),
  2887 => std_logic_vector'(x"00000000"),
  2888 => std_logic_vector'(x"00000000"),
  2889 => std_logic_vector'(x"00000000"),
  2890 => std_logic_vector'(x"00000000"),
  2891 => std_logic_vector'(x"00000000"),
  2892 => std_logic_vector'(x"00000000"),
  2893 => std_logic_vector'(x"00000000"),
  2894 => std_logic_vector'(x"00000000"),
  2895 => std_logic_vector'(x"00000000"),
  2896 => std_logic_vector'(x"00000000"),
  2897 => std_logic_vector'(x"00000000"),
  2898 => std_logic_vector'(x"00000000"),
  2899 => std_logic_vector'(x"00000000"),
  2900 => std_logic_vector'(x"00000000"),
  2901 => std_logic_vector'(x"00000000"),
  2902 => std_logic_vector'(x"00000000"),
  2903 => std_logic_vector'(x"00000000"),
  2904 => std_logic_vector'(x"00000000"),
  2905 => std_logic_vector'(x"00000000"),
  2906 => std_logic_vector'(x"00000000"),
  2907 => std_logic_vector'(x"00000000"),
  2908 => std_logic_vector'(x"00000000"),
  2909 => std_logic_vector'(x"00000000"),
  2910 => std_logic_vector'(x"00000000"),
  2911 => std_logic_vector'(x"00000000"),
  2912 => std_logic_vector'(x"00000000"),
  2913 => std_logic_vector'(x"00000000"),
  2914 => std_logic_vector'(x"00000000"),
  2915 => std_logic_vector'(x"00000000"),
  2916 => std_logic_vector'(x"00000000"),
  2917 => std_logic_vector'(x"00000000"),
  2918 => std_logic_vector'(x"00000000"),
  2919 => std_logic_vector'(x"00000000"),
  2920 => std_logic_vector'(x"00000000"),
  2921 => std_logic_vector'(x"00000000"),
  2922 => std_logic_vector'(x"00000000"),
  2923 => std_logic_vector'(x"00000000"),
  2924 => std_logic_vector'(x"00000000"),
  2925 => std_logic_vector'(x"00000000"),
  2926 => std_logic_vector'(x"00000000"),
  2927 => std_logic_vector'(x"00000000"),
  2928 => std_logic_vector'(x"00000000"),
  2929 => std_logic_vector'(x"00000000"),
  2930 => std_logic_vector'(x"00000000"),
  2931 => std_logic_vector'(x"00000000"),
  2932 => std_logic_vector'(x"00000000"),
  2933 => std_logic_vector'(x"00000000"),
  2934 => std_logic_vector'(x"00000000"),
  2935 => std_logic_vector'(x"00000000"),
  2936 => std_logic_vector'(x"00000000"),
  2937 => std_logic_vector'(x"00000000"),
  2938 => std_logic_vector'(x"00000000"),
  2939 => std_logic_vector'(x"00000000"),
  2940 => std_logic_vector'(x"00000000"),
  2941 => std_logic_vector'(x"00000000"),
  2942 => std_logic_vector'(x"00000000"),
  2943 => std_logic_vector'(x"00000000"),
  2944 => std_logic_vector'(x"00000000"),
  2945 => std_logic_vector'(x"00000000"),
  2946 => std_logic_vector'(x"00000000"),
  2947 => std_logic_vector'(x"00000000"),
  2948 => std_logic_vector'(x"00000000"),
  2949 => std_logic_vector'(x"00000000"),
  2950 => std_logic_vector'(x"00000000"),
  2951 => std_logic_vector'(x"00000000"),
  2952 => std_logic_vector'(x"00000000"),
  2953 => std_logic_vector'(x"00000000"),
  2954 => std_logic_vector'(x"00000000"),
  2955 => std_logic_vector'(x"00000000"),
  2956 => std_logic_vector'(x"00000000"),
  2957 => std_logic_vector'(x"00000000"),
  2958 => std_logic_vector'(x"00000000"),
  2959 => std_logic_vector'(x"00000000"),
  2960 => std_logic_vector'(x"00000000"),
  2961 => std_logic_vector'(x"00000000"),
  2962 => std_logic_vector'(x"00000000"),
  2963 => std_logic_vector'(x"00000000"),
  2964 => std_logic_vector'(x"00000000"),
  2965 => std_logic_vector'(x"00000000"),
  2966 => std_logic_vector'(x"00000000"),
  2967 => std_logic_vector'(x"00000000"),
  2968 => std_logic_vector'(x"00000000"),
  2969 => std_logic_vector'(x"00000000"),
  2970 => std_logic_vector'(x"00000000"),
  2971 => std_logic_vector'(x"00000000"),
  2972 => std_logic_vector'(x"00000000"),
  2973 => std_logic_vector'(x"00000000"),
  2974 => std_logic_vector'(x"00000000"),
  2975 => std_logic_vector'(x"00000000"),
  2976 => std_logic_vector'(x"00000000"),
  2977 => std_logic_vector'(x"00000000"),
  2978 => std_logic_vector'(x"00000000"),
  2979 => std_logic_vector'(x"00000000"),
  2980 => std_logic_vector'(x"00000000"),
  2981 => std_logic_vector'(x"00000000"),
  2982 => std_logic_vector'(x"00000000"),
  2983 => std_logic_vector'(x"00000000"),
  2984 => std_logic_vector'(x"00000000"),
  2985 => std_logic_vector'(x"00000000"),
  2986 => std_logic_vector'(x"00000000"),
  2987 => std_logic_vector'(x"00000000"),
  2988 => std_logic_vector'(x"00000000"),
  2989 => std_logic_vector'(x"00000000"),
  2990 => std_logic_vector'(x"00000000"),
  2991 => std_logic_vector'(x"00000000"),
  2992 => std_logic_vector'(x"00000000"),
  2993 => std_logic_vector'(x"00000000"),
  2994 => std_logic_vector'(x"00000000"),
  2995 => std_logic_vector'(x"00000000"),
  2996 => std_logic_vector'(x"00000000"),
  2997 => std_logic_vector'(x"00000000"),
  2998 => std_logic_vector'(x"00000000"),
  2999 => std_logic_vector'(x"00000000"),
  3000 => std_logic_vector'(x"00000000"),
  3001 => std_logic_vector'(x"00000000"),
  3002 => std_logic_vector'(x"00000000"),
  3003 => std_logic_vector'(x"00000000"),
  3004 => std_logic_vector'(x"00000000"),
  3005 => std_logic_vector'(x"00000000"),
  3006 => std_logic_vector'(x"00000000"),
  3007 => std_logic_vector'(x"00000000"),
  3008 => std_logic_vector'(x"00000000"),
  3009 => std_logic_vector'(x"00000000"),
  3010 => std_logic_vector'(x"00000000"),
  3011 => std_logic_vector'(x"00000000"),
  3012 => std_logic_vector'(x"00000000"),
  3013 => std_logic_vector'(x"00000000"),
  3014 => std_logic_vector'(x"00000000"),
  3015 => std_logic_vector'(x"00000000"),
  3016 => std_logic_vector'(x"00000000"),
  3017 => std_logic_vector'(x"00000000"),
  3018 => std_logic_vector'(x"00000000"),
  3019 => std_logic_vector'(x"00000000"),
  3020 => std_logic_vector'(x"00000000"),
  3021 => std_logic_vector'(x"00000000"),
  3022 => std_logic_vector'(x"00000000"),
  3023 => std_logic_vector'(x"00000000"),
  3024 => std_logic_vector'(x"00000000"),
  3025 => std_logic_vector'(x"00000000"),
  3026 => std_logic_vector'(x"00000000"),
  3027 => std_logic_vector'(x"00000000"),
  3028 => std_logic_vector'(x"00000000"),
  3029 => std_logic_vector'(x"00000000"),
  3030 => std_logic_vector'(x"00000000"),
  3031 => std_logic_vector'(x"00000000"),
  3032 => std_logic_vector'(x"00000000"),
  3033 => std_logic_vector'(x"00000000"),
  3034 => std_logic_vector'(x"00000000"),
  3035 => std_logic_vector'(x"00000000"),
  3036 => std_logic_vector'(x"00000000"),
  3037 => std_logic_vector'(x"00000000"),
  3038 => std_logic_vector'(x"00000000"),
  3039 => std_logic_vector'(x"00000000"),
  3040 => std_logic_vector'(x"00000000"),
  3041 => std_logic_vector'(x"00000000"),
  3042 => std_logic_vector'(x"00000000"),
  3043 => std_logic_vector'(x"00000000"),
  3044 => std_logic_vector'(x"00000000"),
  3045 => std_logic_vector'(x"00000000"),
  3046 => std_logic_vector'(x"00000000"),
  3047 => std_logic_vector'(x"00000000"),
  3048 => std_logic_vector'(x"00000000"),
  3049 => std_logic_vector'(x"00000000"),
  3050 => std_logic_vector'(x"00000000"),
  3051 => std_logic_vector'(x"00000000"),
  3052 => std_logic_vector'(x"00000000"),
  3053 => std_logic_vector'(x"00000000"),
  3054 => std_logic_vector'(x"00000000"),
  3055 => std_logic_vector'(x"00000000"),
  3056 => std_logic_vector'(x"00000000"),
  3057 => std_logic_vector'(x"00000000"),
  3058 => std_logic_vector'(x"00000000"),
  3059 => std_logic_vector'(x"00000000"),
  3060 => std_logic_vector'(x"00000000"),
  3061 => std_logic_vector'(x"00000000"),
  3062 => std_logic_vector'(x"00000000"),
  3063 => std_logic_vector'(x"00000000"),
  3064 => std_logic_vector'(x"00000000"),
  3065 => std_logic_vector'(x"00000000"),
  3066 => std_logic_vector'(x"00000000"),
  3067 => std_logic_vector'(x"00000000"),
  3068 => std_logic_vector'(x"00000000"),
  3069 => std_logic_vector'(x"00000000"),
  3070 => std_logic_vector'(x"00000000"),
  3071 => std_logic_vector'(x"00000000"),
  3072 => std_logic_vector'(x"00000000"),
  3073 => std_logic_vector'(x"00000000"),
  3074 => std_logic_vector'(x"00000000"),
  3075 => std_logic_vector'(x"00000000"),
  3076 => std_logic_vector'(x"00000000"),
  3077 => std_logic_vector'(x"00000000"),
  3078 => std_logic_vector'(x"00000000"),
  3079 => std_logic_vector'(x"00000000"),
  3080 => std_logic_vector'(x"00000000"),
  3081 => std_logic_vector'(x"00000000"),
  3082 => std_logic_vector'(x"00000000"),
  3083 => std_logic_vector'(x"00000000"),
  3084 => std_logic_vector'(x"00000000"),
  3085 => std_logic_vector'(x"00000000"),
  3086 => std_logic_vector'(x"00000000"),
  3087 => std_logic_vector'(x"00000000"),
  3088 => std_logic_vector'(x"00000000"),
  3089 => std_logic_vector'(x"00000000"),
  3090 => std_logic_vector'(x"00000000"),
  3091 => std_logic_vector'(x"00000000"),
  3092 => std_logic_vector'(x"00000000"),
  3093 => std_logic_vector'(x"00000000"),
  3094 => std_logic_vector'(x"00000000"),
  3095 => std_logic_vector'(x"00000000"),
  3096 => std_logic_vector'(x"00000000"),
  3097 => std_logic_vector'(x"00000000"),
  3098 => std_logic_vector'(x"00000000"),
  3099 => std_logic_vector'(x"00000000"),
  3100 => std_logic_vector'(x"00000000"),
  3101 => std_logic_vector'(x"00000000"),
  3102 => std_logic_vector'(x"00000000"),
  3103 => std_logic_vector'(x"00000000"),
  3104 => std_logic_vector'(x"00000000"),
  3105 => std_logic_vector'(x"00000000"),
  3106 => std_logic_vector'(x"00000000"),
  3107 => std_logic_vector'(x"00000000"),
  3108 => std_logic_vector'(x"00000000"),
  3109 => std_logic_vector'(x"00000000"),
  3110 => std_logic_vector'(x"00000000"),
  3111 => std_logic_vector'(x"00000000"),
  3112 => std_logic_vector'(x"00000000"),
  3113 => std_logic_vector'(x"00000000"),
  3114 => std_logic_vector'(x"00000000"),
  3115 => std_logic_vector'(x"00000000"),
  3116 => std_logic_vector'(x"00000000"),
  3117 => std_logic_vector'(x"00000000"),
  3118 => std_logic_vector'(x"00000000"),
  3119 => std_logic_vector'(x"00000000"),
  3120 => std_logic_vector'(x"00000000"),
  3121 => std_logic_vector'(x"00000000"),
  3122 => std_logic_vector'(x"00000000"),
  3123 => std_logic_vector'(x"00000000"),
  3124 => std_logic_vector'(x"00000000"),
  3125 => std_logic_vector'(x"00000000"),
  3126 => std_logic_vector'(x"00000000"),
  3127 => std_logic_vector'(x"00000000"),
  3128 => std_logic_vector'(x"00000000"),
  3129 => std_logic_vector'(x"00000000"),
  3130 => std_logic_vector'(x"00000000"),
  3131 => std_logic_vector'(x"00000000"),
  3132 => std_logic_vector'(x"00000000"),
  3133 => std_logic_vector'(x"00000000"),
  3134 => std_logic_vector'(x"00000000"),
  3135 => std_logic_vector'(x"00000000"),
  3136 => std_logic_vector'(x"00000000"),
  3137 => std_logic_vector'(x"00000000"),
  3138 => std_logic_vector'(x"00000000"),
  3139 => std_logic_vector'(x"00000000"),
  3140 => std_logic_vector'(x"00000000"),
  3141 => std_logic_vector'(x"00000000"),
  3142 => std_logic_vector'(x"00000000"),
  3143 => std_logic_vector'(x"00000000"),
  3144 => std_logic_vector'(x"00000000"),
  3145 => std_logic_vector'(x"00000000"),
  3146 => std_logic_vector'(x"00000000"),
  3147 => std_logic_vector'(x"00000000"),
  3148 => std_logic_vector'(x"00000000"),
  3149 => std_logic_vector'(x"00000000"),
  3150 => std_logic_vector'(x"00000000"),
  3151 => std_logic_vector'(x"00000000"),
  3152 => std_logic_vector'(x"00000000"),
  3153 => std_logic_vector'(x"00000000"),
  3154 => std_logic_vector'(x"00000000"),
  3155 => std_logic_vector'(x"00000000"),
  3156 => std_logic_vector'(x"00000000"),
  3157 => std_logic_vector'(x"00000000"),
  3158 => std_logic_vector'(x"00000000"),
  3159 => std_logic_vector'(x"00000000"),
  3160 => std_logic_vector'(x"00000000"),
  3161 => std_logic_vector'(x"00000000"),
  3162 => std_logic_vector'(x"00000000"),
  3163 => std_logic_vector'(x"00000000"),
  3164 => std_logic_vector'(x"00000000"),
  3165 => std_logic_vector'(x"00000000"),
  3166 => std_logic_vector'(x"00000000"),
  3167 => std_logic_vector'(x"00000000"),
  3168 => std_logic_vector'(x"00000000"),
  3169 => std_logic_vector'(x"00000000"),
  3170 => std_logic_vector'(x"00000000"),
  3171 => std_logic_vector'(x"00000000"),
  3172 => std_logic_vector'(x"00000000"),
  3173 => std_logic_vector'(x"00000000"),
  3174 => std_logic_vector'(x"00000000"),
  3175 => std_logic_vector'(x"00000000"),
  3176 => std_logic_vector'(x"00000000"),
  3177 => std_logic_vector'(x"00000000"),
  3178 => std_logic_vector'(x"00000000"),
  3179 => std_logic_vector'(x"00000000"),
  3180 => std_logic_vector'(x"00000000"),
  3181 => std_logic_vector'(x"00000000"),
  3182 => std_logic_vector'(x"00000000"),
  3183 => std_logic_vector'(x"00000000"),
  3184 => std_logic_vector'(x"00000000"),
  3185 => std_logic_vector'(x"00000000"),
  3186 => std_logic_vector'(x"00000000"),
  3187 => std_logic_vector'(x"00000000"),
  3188 => std_logic_vector'(x"00000000"),
  3189 => std_logic_vector'(x"00000000"),
  3190 => std_logic_vector'(x"00000000"),
  3191 => std_logic_vector'(x"00000000"),
  3192 => std_logic_vector'(x"00000000"),
  3193 => std_logic_vector'(x"00000000"),
  3194 => std_logic_vector'(x"00000000"),
  3195 => std_logic_vector'(x"00000000"),
  3196 => std_logic_vector'(x"00000000"),
  3197 => std_logic_vector'(x"00000000"),
  3198 => std_logic_vector'(x"00000000"),
  3199 => std_logic_vector'(x"00000000"),
  3200 => std_logic_vector'(x"00000000"),
  3201 => std_logic_vector'(x"00000000"),
  3202 => std_logic_vector'(x"00000000"),
  3203 => std_logic_vector'(x"00000000"),
  3204 => std_logic_vector'(x"00000000"),
  3205 => std_logic_vector'(x"00000000"),
  3206 => std_logic_vector'(x"00000000"),
  3207 => std_logic_vector'(x"00000000"),
  3208 => std_logic_vector'(x"00000000"),
  3209 => std_logic_vector'(x"00000000"),
  3210 => std_logic_vector'(x"00000000"),
  3211 => std_logic_vector'(x"00000000"),
  3212 => std_logic_vector'(x"00000000"),
  3213 => std_logic_vector'(x"00000000"),
  3214 => std_logic_vector'(x"00000000"),
  3215 => std_logic_vector'(x"00000000"),
  3216 => std_logic_vector'(x"00000000"),
  3217 => std_logic_vector'(x"00000000"),
  3218 => std_logic_vector'(x"00000000"),
  3219 => std_logic_vector'(x"00000000"),
  3220 => std_logic_vector'(x"00000000"),
  3221 => std_logic_vector'(x"00000000"),
  3222 => std_logic_vector'(x"00000000"),
  3223 => std_logic_vector'(x"00000000"),
  3224 => std_logic_vector'(x"00000000"),
  3225 => std_logic_vector'(x"00000000"),
  3226 => std_logic_vector'(x"00000000"),
  3227 => std_logic_vector'(x"00000000"),
  3228 => std_logic_vector'(x"00000000"),
  3229 => std_logic_vector'(x"00000000"),
  3230 => std_logic_vector'(x"00000000"),
  3231 => std_logic_vector'(x"00000000"),
  3232 => std_logic_vector'(x"00000000"),
  3233 => std_logic_vector'(x"00000000"),
  3234 => std_logic_vector'(x"00000000"),
  3235 => std_logic_vector'(x"00000000"),
  3236 => std_logic_vector'(x"00000000"),
  3237 => std_logic_vector'(x"00000000"),
  3238 => std_logic_vector'(x"00000000"),
  3239 => std_logic_vector'(x"00000000"),
  3240 => std_logic_vector'(x"00000000"),
  3241 => std_logic_vector'(x"00000000"),
  3242 => std_logic_vector'(x"00000000"),
  3243 => std_logic_vector'(x"00000000"),
  3244 => std_logic_vector'(x"00000000"),
  3245 => std_logic_vector'(x"00000000"),
  3246 => std_logic_vector'(x"00000000"),
  3247 => std_logic_vector'(x"00000000"),
  3248 => std_logic_vector'(x"00000000"),
  3249 => std_logic_vector'(x"00000000"),
  3250 => std_logic_vector'(x"00000000"),
  3251 => std_logic_vector'(x"00000000"),
  3252 => std_logic_vector'(x"00000000"),
  3253 => std_logic_vector'(x"00000000"),
  3254 => std_logic_vector'(x"00000000"),
  3255 => std_logic_vector'(x"00000000"),
  3256 => std_logic_vector'(x"00000000"),
  3257 => std_logic_vector'(x"00000000"),
  3258 => std_logic_vector'(x"00000000"),
  3259 => std_logic_vector'(x"00000000"),
  3260 => std_logic_vector'(x"00000000"),
  3261 => std_logic_vector'(x"00000000"),
  3262 => std_logic_vector'(x"00000000"),
  3263 => std_logic_vector'(x"00000000"),
  3264 => std_logic_vector'(x"00000000"),
  3265 => std_logic_vector'(x"00000000"),
  3266 => std_logic_vector'(x"00000000"),
  3267 => std_logic_vector'(x"00000000"),
  3268 => std_logic_vector'(x"00000000"),
  3269 => std_logic_vector'(x"00000000"),
  3270 => std_logic_vector'(x"00000000"),
  3271 => std_logic_vector'(x"00000000"),
  3272 => std_logic_vector'(x"00000000"),
  3273 => std_logic_vector'(x"00000000"),
  3274 => std_logic_vector'(x"00000000"),
  3275 => std_logic_vector'(x"00000000"),
  3276 => std_logic_vector'(x"00000000"),
  3277 => std_logic_vector'(x"00000000"),
  3278 => std_logic_vector'(x"00000000"),
  3279 => std_logic_vector'(x"00000000"),
  3280 => std_logic_vector'(x"00000000"),
  3281 => std_logic_vector'(x"00000000"),
  3282 => std_logic_vector'(x"00000000"),
  3283 => std_logic_vector'(x"00000000"),
  3284 => std_logic_vector'(x"00000000"),
  3285 => std_logic_vector'(x"00000000"),
  3286 => std_logic_vector'(x"00000000"),
  3287 => std_logic_vector'(x"00000000"),
  3288 => std_logic_vector'(x"00000000"),
  3289 => std_logic_vector'(x"00000000"),
  3290 => std_logic_vector'(x"00000000"),
  3291 => std_logic_vector'(x"00000000"),
  3292 => std_logic_vector'(x"00000000"),
  3293 => std_logic_vector'(x"00000000"),
  3294 => std_logic_vector'(x"00000000"),
  3295 => std_logic_vector'(x"00000000"),
  3296 => std_logic_vector'(x"00000000"),
  3297 => std_logic_vector'(x"00000000"),
  3298 => std_logic_vector'(x"00000000"),
  3299 => std_logic_vector'(x"00000000"),
  3300 => std_logic_vector'(x"00000000"),
  3301 => std_logic_vector'(x"00000000"),
  3302 => std_logic_vector'(x"00000000"),
  3303 => std_logic_vector'(x"00000000"),
  3304 => std_logic_vector'(x"00000000"),
  3305 => std_logic_vector'(x"00000000"),
  3306 => std_logic_vector'(x"00000000"),
  3307 => std_logic_vector'(x"00000000"),
  3308 => std_logic_vector'(x"00000000"),
  3309 => std_logic_vector'(x"00000000"),
  3310 => std_logic_vector'(x"00000000"),
  3311 => std_logic_vector'(x"00000000"),
  3312 => std_logic_vector'(x"00000000"),
  3313 => std_logic_vector'(x"00000000"),
  3314 => std_logic_vector'(x"00000000"),
  3315 => std_logic_vector'(x"00000000"),
  3316 => std_logic_vector'(x"00000000"),
  3317 => std_logic_vector'(x"00000000"),
  3318 => std_logic_vector'(x"00000000"),
  3319 => std_logic_vector'(x"00000000"),
  3320 => std_logic_vector'(x"00000000"),
  3321 => std_logic_vector'(x"00000000"),
  3322 => std_logic_vector'(x"00000000"),
  3323 => std_logic_vector'(x"00000000"),
  3324 => std_logic_vector'(x"00000000"),
  3325 => std_logic_vector'(x"00000000"),
  3326 => std_logic_vector'(x"00000000"),
  3327 => std_logic_vector'(x"00000000"),
  3328 => std_logic_vector'(x"00000000"),
  3329 => std_logic_vector'(x"00000000"),
  3330 => std_logic_vector'(x"00000000"),
  3331 => std_logic_vector'(x"00000000"),
  3332 => std_logic_vector'(x"00000000"),
  3333 => std_logic_vector'(x"00000000"),
  3334 => std_logic_vector'(x"00000000"),
  3335 => std_logic_vector'(x"00000000"),
  3336 => std_logic_vector'(x"00000000"),
  3337 => std_logic_vector'(x"00000000"),
  3338 => std_logic_vector'(x"00000000"),
  3339 => std_logic_vector'(x"00000000"),
  3340 => std_logic_vector'(x"00000000"),
  3341 => std_logic_vector'(x"00000000"),
  3342 => std_logic_vector'(x"00000000"),
  3343 => std_logic_vector'(x"00000000"),
  3344 => std_logic_vector'(x"00000000"),
  3345 => std_logic_vector'(x"00000000"),
  3346 => std_logic_vector'(x"00000000"),
  3347 => std_logic_vector'(x"00000000"),
  3348 => std_logic_vector'(x"00000000"),
  3349 => std_logic_vector'(x"00000000"),
  3350 => std_logic_vector'(x"00000000"),
  3351 => std_logic_vector'(x"00000000"),
  3352 => std_logic_vector'(x"00000000"),
  3353 => std_logic_vector'(x"00000000"),
  3354 => std_logic_vector'(x"00000000"),
  3355 => std_logic_vector'(x"00000000"),
  3356 => std_logic_vector'(x"00000000"),
  3357 => std_logic_vector'(x"00000000"),
  3358 => std_logic_vector'(x"00000000"),
  3359 => std_logic_vector'(x"00000000"),
  3360 => std_logic_vector'(x"00000000"),
  3361 => std_logic_vector'(x"00000000"),
  3362 => std_logic_vector'(x"00000000"),
  3363 => std_logic_vector'(x"00000000"),
  3364 => std_logic_vector'(x"00000000"),
  3365 => std_logic_vector'(x"00000000"),
  3366 => std_logic_vector'(x"00000000"),
  3367 => std_logic_vector'(x"00000000"),
  3368 => std_logic_vector'(x"00000000"),
  3369 => std_logic_vector'(x"00000000"),
  3370 => std_logic_vector'(x"00000000"),
  3371 => std_logic_vector'(x"00000000"),
  3372 => std_logic_vector'(x"00000000"),
  3373 => std_logic_vector'(x"00000000"),
  3374 => std_logic_vector'(x"00000000"),
  3375 => std_logic_vector'(x"00000000"),
  3376 => std_logic_vector'(x"00000000"),
  3377 => std_logic_vector'(x"00000000"),
  3378 => std_logic_vector'(x"00000000"),
  3379 => std_logic_vector'(x"00000000"),
  3380 => std_logic_vector'(x"00000000"),
  3381 => std_logic_vector'(x"00000000"),
  3382 => std_logic_vector'(x"00000000"),
  3383 => std_logic_vector'(x"00000000"),
  3384 => std_logic_vector'(x"00000000"),
  3385 => std_logic_vector'(x"00000000"),
  3386 => std_logic_vector'(x"00000000"),
  3387 => std_logic_vector'(x"00000000"),
  3388 => std_logic_vector'(x"00000000"),
  3389 => std_logic_vector'(x"00000000"),
  3390 => std_logic_vector'(x"00000000"),
  3391 => std_logic_vector'(x"00000000"),
  3392 => std_logic_vector'(x"00000000"),
  3393 => std_logic_vector'(x"00000000"),
  3394 => std_logic_vector'(x"00000000"),
  3395 => std_logic_vector'(x"00000000"),
  3396 => std_logic_vector'(x"00000000"),
  3397 => std_logic_vector'(x"00000000"),
  3398 => std_logic_vector'(x"00000000"),
  3399 => std_logic_vector'(x"00000000"),
  3400 => std_logic_vector'(x"00000000"),
  3401 => std_logic_vector'(x"00000000"),
  3402 => std_logic_vector'(x"00000000"),
  3403 => std_logic_vector'(x"00000000"),
  3404 => std_logic_vector'(x"00000000"),
  3405 => std_logic_vector'(x"00000000"),
  3406 => std_logic_vector'(x"00000000"),
  3407 => std_logic_vector'(x"00000000"),
  3408 => std_logic_vector'(x"00000000"),
  3409 => std_logic_vector'(x"00000000"),
  3410 => std_logic_vector'(x"00000000"),
  3411 => std_logic_vector'(x"00000000"),
  3412 => std_logic_vector'(x"00000000"),
  3413 => std_logic_vector'(x"00000000"),
  3414 => std_logic_vector'(x"00000000"),
  3415 => std_logic_vector'(x"00000000"),
  3416 => std_logic_vector'(x"00000000"),
  3417 => std_logic_vector'(x"00000000"),
  3418 => std_logic_vector'(x"00000000"),
  3419 => std_logic_vector'(x"00000000"),
  3420 => std_logic_vector'(x"00000000"),
  3421 => std_logic_vector'(x"00000000"),
  3422 => std_logic_vector'(x"00000000"),
  3423 => std_logic_vector'(x"00000000"),
  3424 => std_logic_vector'(x"00000000"),
  3425 => std_logic_vector'(x"00000000"),
  3426 => std_logic_vector'(x"00000000"),
  3427 => std_logic_vector'(x"00000000"),
  3428 => std_logic_vector'(x"00000000"),
  3429 => std_logic_vector'(x"00000000"),
  3430 => std_logic_vector'(x"00000000"),
  3431 => std_logic_vector'(x"00000000"),
  3432 => std_logic_vector'(x"00000000"),
  3433 => std_logic_vector'(x"00000000"),
  3434 => std_logic_vector'(x"00000000"),
  3435 => std_logic_vector'(x"00000000"),
  3436 => std_logic_vector'(x"00000000"),
  3437 => std_logic_vector'(x"00000000"),
  3438 => std_logic_vector'(x"00000000"),
  3439 => std_logic_vector'(x"00000000"),
  3440 => std_logic_vector'(x"00000000"),
  3441 => std_logic_vector'(x"00000000"),
  3442 => std_logic_vector'(x"00000000"),
  3443 => std_logic_vector'(x"00000000"),
  3444 => std_logic_vector'(x"00000000"),
  3445 => std_logic_vector'(x"00000000"),
  3446 => std_logic_vector'(x"00000000"),
  3447 => std_logic_vector'(x"00000000"),
  3448 => std_logic_vector'(x"00000000"),
  3449 => std_logic_vector'(x"00000000"),
  3450 => std_logic_vector'(x"00000000"),
  3451 => std_logic_vector'(x"00000000"),
  3452 => std_logic_vector'(x"00000000"),
  3453 => std_logic_vector'(x"00000000"),
  3454 => std_logic_vector'(x"00000000"),
  3455 => std_logic_vector'(x"00000000"),
  3456 => std_logic_vector'(x"00000000"),
  3457 => std_logic_vector'(x"00000000"),
  3458 => std_logic_vector'(x"00000000"),
  3459 => std_logic_vector'(x"00000000"),
  3460 => std_logic_vector'(x"00000000"),
  3461 => std_logic_vector'(x"00000000"),
  3462 => std_logic_vector'(x"00000000"),
  3463 => std_logic_vector'(x"00000000"),
  3464 => std_logic_vector'(x"00000000"),
  3465 => std_logic_vector'(x"00000000"),
  3466 => std_logic_vector'(x"00000000"),
  3467 => std_logic_vector'(x"00000000"),
  3468 => std_logic_vector'(x"00000000"),
  3469 => std_logic_vector'(x"00000000"),
  3470 => std_logic_vector'(x"00000000"),
  3471 => std_logic_vector'(x"00000000"),
  3472 => std_logic_vector'(x"00000000"),
  3473 => std_logic_vector'(x"00000000"),
  3474 => std_logic_vector'(x"00000000"),
  3475 => std_logic_vector'(x"00000000"),
  3476 => std_logic_vector'(x"00000000"),
  3477 => std_logic_vector'(x"00000000"),
  3478 => std_logic_vector'(x"00000000"),
  3479 => std_logic_vector'(x"00000000"),
  3480 => std_logic_vector'(x"00000000"),
  3481 => std_logic_vector'(x"00000000"),
  3482 => std_logic_vector'(x"00000000"),
  3483 => std_logic_vector'(x"00000000"),
  3484 => std_logic_vector'(x"00000000"),
  3485 => std_logic_vector'(x"00000000"),
  3486 => std_logic_vector'(x"00000000"),
  3487 => std_logic_vector'(x"00000000"),
  3488 => std_logic_vector'(x"00000000"),
  3489 => std_logic_vector'(x"00000000"),
  3490 => std_logic_vector'(x"00000000"),
  3491 => std_logic_vector'(x"00000000"),
  3492 => std_logic_vector'(x"00000000"),
  3493 => std_logic_vector'(x"00000000"),
  3494 => std_logic_vector'(x"00000000"),
  3495 => std_logic_vector'(x"00000000"),
  3496 => std_logic_vector'(x"00000000"),
  3497 => std_logic_vector'(x"00000000"),
  3498 => std_logic_vector'(x"00000000"),
  3499 => std_logic_vector'(x"00000000"),
  3500 => std_logic_vector'(x"00000000"),
  3501 => std_logic_vector'(x"00000000"),
  3502 => std_logic_vector'(x"00000000"),
  3503 => std_logic_vector'(x"00000000"),
  3504 => std_logic_vector'(x"00000000"),
  3505 => std_logic_vector'(x"00000000"),
  3506 => std_logic_vector'(x"00000000"),
  3507 => std_logic_vector'(x"00000000"),
  3508 => std_logic_vector'(x"00000000"),
  3509 => std_logic_vector'(x"00000000"),
  3510 => std_logic_vector'(x"00000000"),
  3511 => std_logic_vector'(x"00000000"),
  3512 => std_logic_vector'(x"00000000"),
  3513 => std_logic_vector'(x"00000000"),
  3514 => std_logic_vector'(x"00000000"),
  3515 => std_logic_vector'(x"00000000"),
  3516 => std_logic_vector'(x"00000000"),
  3517 => std_logic_vector'(x"00000000"),
  3518 => std_logic_vector'(x"00000000"),
  3519 => std_logic_vector'(x"00000000"),
  3520 => std_logic_vector'(x"00000000"),
  3521 => std_logic_vector'(x"00000000"),
  3522 => std_logic_vector'(x"00000000"),
  3523 => std_logic_vector'(x"00000000"),
  3524 => std_logic_vector'(x"00000000"),
  3525 => std_logic_vector'(x"00000000"),
  3526 => std_logic_vector'(x"00000000"),
  3527 => std_logic_vector'(x"00000000"),
  3528 => std_logic_vector'(x"00000000"),
  3529 => std_logic_vector'(x"00000000"),
  3530 => std_logic_vector'(x"00000000"),
  3531 => std_logic_vector'(x"00000000"),
  3532 => std_logic_vector'(x"00000000"),
  3533 => std_logic_vector'(x"00000000"),
  3534 => std_logic_vector'(x"00000000"),
  3535 => std_logic_vector'(x"00000000"),
  3536 => std_logic_vector'(x"00000000"),
  3537 => std_logic_vector'(x"00000000"),
  3538 => std_logic_vector'(x"00000000"),
  3539 => std_logic_vector'(x"00000000"),
  3540 => std_logic_vector'(x"00000000"),
  3541 => std_logic_vector'(x"00000000"),
  3542 => std_logic_vector'(x"00000000"),
  3543 => std_logic_vector'(x"00000000"),
  3544 => std_logic_vector'(x"00000000"),
  3545 => std_logic_vector'(x"00000000"),
  3546 => std_logic_vector'(x"00000000"),
  3547 => std_logic_vector'(x"00000000"),
  3548 => std_logic_vector'(x"00000000"),
  3549 => std_logic_vector'(x"00000000"),
  3550 => std_logic_vector'(x"00000000"),
  3551 => std_logic_vector'(x"00000000"),
  3552 => std_logic_vector'(x"00000000"),
  3553 => std_logic_vector'(x"00000000"),
  3554 => std_logic_vector'(x"00000000"),
  3555 => std_logic_vector'(x"00000000"),
  3556 => std_logic_vector'(x"00000000"),
  3557 => std_logic_vector'(x"00000000"),
  3558 => std_logic_vector'(x"00000000"),
  3559 => std_logic_vector'(x"00000000"),
  3560 => std_logic_vector'(x"00000000"),
  3561 => std_logic_vector'(x"00000000"),
  3562 => std_logic_vector'(x"00000000"),
  3563 => std_logic_vector'(x"00000000"),
  3564 => std_logic_vector'(x"00000000"),
  3565 => std_logic_vector'(x"00000000"),
  3566 => std_logic_vector'(x"00000000"),
  3567 => std_logic_vector'(x"00000000"),
  3568 => std_logic_vector'(x"00000000"),
  3569 => std_logic_vector'(x"00000000"),
  3570 => std_logic_vector'(x"00000000"),
  3571 => std_logic_vector'(x"00000000"),
  3572 => std_logic_vector'(x"00000000"),
  3573 => std_logic_vector'(x"00000000"),
  3574 => std_logic_vector'(x"00000000"),
  3575 => std_logic_vector'(x"00000000"),
  3576 => std_logic_vector'(x"00000000"),
  3577 => std_logic_vector'(x"00000000"),
  3578 => std_logic_vector'(x"00000000"),
  3579 => std_logic_vector'(x"00000000"),
  3580 => std_logic_vector'(x"00000000"),
  3581 => std_logic_vector'(x"00000000"),
  3582 => std_logic_vector'(x"00000000"),
  3583 => std_logic_vector'(x"00000000"),
  3584 => std_logic_vector'(x"00000000"),
  3585 => std_logic_vector'(x"00000000"),
  3586 => std_logic_vector'(x"00000000"),
  3587 => std_logic_vector'(x"00000000"),
  3588 => std_logic_vector'(x"00000000"),
  3589 => std_logic_vector'(x"00000000"),
  3590 => std_logic_vector'(x"00000000"),
  3591 => std_logic_vector'(x"00000000"),
  3592 => std_logic_vector'(x"00000000"),
  3593 => std_logic_vector'(x"00000000"),
  3594 => std_logic_vector'(x"00000000"),
  3595 => std_logic_vector'(x"00000000"),
  3596 => std_logic_vector'(x"00000000"),
  3597 => std_logic_vector'(x"00000000"),
  3598 => std_logic_vector'(x"00000000"),
  3599 => std_logic_vector'(x"00000000"),
  3600 => std_logic_vector'(x"00000000"),
  3601 => std_logic_vector'(x"00000000"),
  3602 => std_logic_vector'(x"00000000"),
  3603 => std_logic_vector'(x"00000000"),
  3604 => std_logic_vector'(x"00000000"),
  3605 => std_logic_vector'(x"00000000"),
  3606 => std_logic_vector'(x"00000000"),
  3607 => std_logic_vector'(x"00000000"),
  3608 => std_logic_vector'(x"00000000"),
  3609 => std_logic_vector'(x"00000000"),
  3610 => std_logic_vector'(x"00000000"),
  3611 => std_logic_vector'(x"00000000"),
  3612 => std_logic_vector'(x"00000000"),
  3613 => std_logic_vector'(x"00000000"),
  3614 => std_logic_vector'(x"00000000"),
  3615 => std_logic_vector'(x"00000000"),
  3616 => std_logic_vector'(x"00000000"),
  3617 => std_logic_vector'(x"00000000"),
  3618 => std_logic_vector'(x"00000000"),
  3619 => std_logic_vector'(x"00000000"),
  3620 => std_logic_vector'(x"00000000"),
  3621 => std_logic_vector'(x"00000000"),
  3622 => std_logic_vector'(x"00000000"),
  3623 => std_logic_vector'(x"00000000"),
  3624 => std_logic_vector'(x"00000000"),
  3625 => std_logic_vector'(x"00000000"),
  3626 => std_logic_vector'(x"00000000"),
  3627 => std_logic_vector'(x"00000000"),
  3628 => std_logic_vector'(x"00000000"),
  3629 => std_logic_vector'(x"00000000"),
  3630 => std_logic_vector'(x"00000000"),
  3631 => std_logic_vector'(x"00000000"),
  3632 => std_logic_vector'(x"00000000"),
  3633 => std_logic_vector'(x"00000000"),
  3634 => std_logic_vector'(x"00000000"),
  3635 => std_logic_vector'(x"00000000"),
  3636 => std_logic_vector'(x"00000000"),
  3637 => std_logic_vector'(x"00000000"),
  3638 => std_logic_vector'(x"00000000"),
  3639 => std_logic_vector'(x"00000000"),
  3640 => std_logic_vector'(x"00000000"),
  3641 => std_logic_vector'(x"00000000"),
  3642 => std_logic_vector'(x"00000000"),
  3643 => std_logic_vector'(x"00000000"),
  3644 => std_logic_vector'(x"00000000"),
  3645 => std_logic_vector'(x"00000000"),
  3646 => std_logic_vector'(x"00000000"),
  3647 => std_logic_vector'(x"00000000"),
  3648 => std_logic_vector'(x"00000000"),
  3649 => std_logic_vector'(x"00000000"),
  3650 => std_logic_vector'(x"00000000"),
  3651 => std_logic_vector'(x"00000000"),
  3652 => std_logic_vector'(x"00000000"),
  3653 => std_logic_vector'(x"00000000"),
  3654 => std_logic_vector'(x"00000000"),
  3655 => std_logic_vector'(x"00000000"),
  3656 => std_logic_vector'(x"00000000"),
  3657 => std_logic_vector'(x"00000000"),
  3658 => std_logic_vector'(x"00000000"),
  3659 => std_logic_vector'(x"00000000"),
  3660 => std_logic_vector'(x"00000000"),
  3661 => std_logic_vector'(x"00000000"),
  3662 => std_logic_vector'(x"00000000"),
  3663 => std_logic_vector'(x"00000000"),
  3664 => std_logic_vector'(x"00000000"),
  3665 => std_logic_vector'(x"00000000"),
  3666 => std_logic_vector'(x"00000000"),
  3667 => std_logic_vector'(x"00000000"),
  3668 => std_logic_vector'(x"00000000"),
  3669 => std_logic_vector'(x"00000000"),
  3670 => std_logic_vector'(x"00000000"),
  3671 => std_logic_vector'(x"00000000"),
  3672 => std_logic_vector'(x"00000000"),
  3673 => std_logic_vector'(x"00000000"),
  3674 => std_logic_vector'(x"00000000"),
  3675 => std_logic_vector'(x"00000000"),
  3676 => std_logic_vector'(x"00000000"),
  3677 => std_logic_vector'(x"00000000"),
  3678 => std_logic_vector'(x"00000000"),
  3679 => std_logic_vector'(x"00000000"),
  3680 => std_logic_vector'(x"00000000"),
  3681 => std_logic_vector'(x"00000000"),
  3682 => std_logic_vector'(x"00000000"),
  3683 => std_logic_vector'(x"00000000"),
  3684 => std_logic_vector'(x"00000000"),
  3685 => std_logic_vector'(x"00000000"),
  3686 => std_logic_vector'(x"00000000"),
  3687 => std_logic_vector'(x"00000000"),
  3688 => std_logic_vector'(x"00000000"),
  3689 => std_logic_vector'(x"00000000"),
  3690 => std_logic_vector'(x"00000000"),
  3691 => std_logic_vector'(x"00000000"),
  3692 => std_logic_vector'(x"00000000"),
  3693 => std_logic_vector'(x"00000000"),
  3694 => std_logic_vector'(x"00000000"),
  3695 => std_logic_vector'(x"00000000"),
  3696 => std_logic_vector'(x"00000000"),
  3697 => std_logic_vector'(x"00000000"),
  3698 => std_logic_vector'(x"00000000"),
  3699 => std_logic_vector'(x"00000000"),
  3700 => std_logic_vector'(x"00000000"),
  3701 => std_logic_vector'(x"00000000"),
  3702 => std_logic_vector'(x"00000000"),
  3703 => std_logic_vector'(x"00000000"),
  3704 => std_logic_vector'(x"00000000"),
  3705 => std_logic_vector'(x"00000000"),
  3706 => std_logic_vector'(x"00000000"),
  3707 => std_logic_vector'(x"00000000"),
  3708 => std_logic_vector'(x"00000000"),
  3709 => std_logic_vector'(x"00000000"),
  3710 => std_logic_vector'(x"00000000"),
  3711 => std_logic_vector'(x"00000000"),
  3712 => std_logic_vector'(x"00000000"),
  3713 => std_logic_vector'(x"00000000"),
  3714 => std_logic_vector'(x"00000000"),
  3715 => std_logic_vector'(x"00000000"),
  3716 => std_logic_vector'(x"00000000"),
  3717 => std_logic_vector'(x"00000000"),
  3718 => std_logic_vector'(x"00000000"),
  3719 => std_logic_vector'(x"00000000"),
  3720 => std_logic_vector'(x"00000000"),
  3721 => std_logic_vector'(x"00000000"),
  3722 => std_logic_vector'(x"00000000"),
  3723 => std_logic_vector'(x"00000000"),
  3724 => std_logic_vector'(x"00000000"),
  3725 => std_logic_vector'(x"00000000"),
  3726 => std_logic_vector'(x"00000000"),
  3727 => std_logic_vector'(x"00000000"),
  3728 => std_logic_vector'(x"00000000"),
  3729 => std_logic_vector'(x"00000000"),
  3730 => std_logic_vector'(x"00000000"),
  3731 => std_logic_vector'(x"00000000"),
  3732 => std_logic_vector'(x"00000000"),
  3733 => std_logic_vector'(x"00000000"),
  3734 => std_logic_vector'(x"00000000"),
  3735 => std_logic_vector'(x"00000000"),
  3736 => std_logic_vector'(x"00000000"),
  3737 => std_logic_vector'(x"00000000"),
  3738 => std_logic_vector'(x"00000000"),
  3739 => std_logic_vector'(x"00000000"),
  3740 => std_logic_vector'(x"00000000"),
  3741 => std_logic_vector'(x"00000000"),
  3742 => std_logic_vector'(x"00000000"),
  3743 => std_logic_vector'(x"00000000"),
  3744 => std_logic_vector'(x"00000000"),
  3745 => std_logic_vector'(x"00000000"),
  3746 => std_logic_vector'(x"00000000"),
  3747 => std_logic_vector'(x"00000000"),
  3748 => std_logic_vector'(x"00000000"),
  3749 => std_logic_vector'(x"00000000"),
  3750 => std_logic_vector'(x"00000000"),
  3751 => std_logic_vector'(x"00000000"),
  3752 => std_logic_vector'(x"00000000"),
  3753 => std_logic_vector'(x"00000000"),
  3754 => std_logic_vector'(x"00000000"),
  3755 => std_logic_vector'(x"00000000"),
  3756 => std_logic_vector'(x"00000000"),
  3757 => std_logic_vector'(x"00000000"),
  3758 => std_logic_vector'(x"00000000"),
  3759 => std_logic_vector'(x"00000000"),
  3760 => std_logic_vector'(x"00000000"),
  3761 => std_logic_vector'(x"00000000"),
  3762 => std_logic_vector'(x"00000000"),
  3763 => std_logic_vector'(x"00000000"),
  3764 => std_logic_vector'(x"00000000"),
  3765 => std_logic_vector'(x"00000000"),
  3766 => std_logic_vector'(x"00000000"),
  3767 => std_logic_vector'(x"00000000"),
  3768 => std_logic_vector'(x"00000000"),
  3769 => std_logic_vector'(x"00000000"),
  3770 => std_logic_vector'(x"00000000"),
  3771 => std_logic_vector'(x"00000000"),
  3772 => std_logic_vector'(x"00000000"),
  3773 => std_logic_vector'(x"00000000"),
  3774 => std_logic_vector'(x"00000000"),
  3775 => std_logic_vector'(x"00000000"),
  3776 => std_logic_vector'(x"00000000"),
  3777 => std_logic_vector'(x"00000000"),
  3778 => std_logic_vector'(x"00000000"),
  3779 => std_logic_vector'(x"00000000"),
  3780 => std_logic_vector'(x"00000000"),
  3781 => std_logic_vector'(x"00000000"),
  3782 => std_logic_vector'(x"00000000"),
  3783 => std_logic_vector'(x"00000000"),
  3784 => std_logic_vector'(x"00000000"),
  3785 => std_logic_vector'(x"00000000"),
  3786 => std_logic_vector'(x"00000000"),
  3787 => std_logic_vector'(x"00000000"),
  3788 => std_logic_vector'(x"00000000"),
  3789 => std_logic_vector'(x"00000000"),
  3790 => std_logic_vector'(x"00000000"),
  3791 => std_logic_vector'(x"00000000"),
  3792 => std_logic_vector'(x"00000000"),
  3793 => std_logic_vector'(x"00000000"),
  3794 => std_logic_vector'(x"00000000"),
  3795 => std_logic_vector'(x"00000000"),
  3796 => std_logic_vector'(x"00000000"),
  3797 => std_logic_vector'(x"00000000"),
  3798 => std_logic_vector'(x"00000000"),
  3799 => std_logic_vector'(x"00000000"),
  3800 => std_logic_vector'(x"00000000"),
  3801 => std_logic_vector'(x"00000000"),
  3802 => std_logic_vector'(x"00000000"),
  3803 => std_logic_vector'(x"00000000"),
  3804 => std_logic_vector'(x"00000000"),
  3805 => std_logic_vector'(x"00000000"),
  3806 => std_logic_vector'(x"00000000"),
  3807 => std_logic_vector'(x"00000000"),
  3808 => std_logic_vector'(x"00000000"),
  3809 => std_logic_vector'(x"00000000"),
  3810 => std_logic_vector'(x"00000000"),
  3811 => std_logic_vector'(x"00000000"),
  3812 => std_logic_vector'(x"00000000"),
  3813 => std_logic_vector'(x"00000000"),
  3814 => std_logic_vector'(x"00000000"),
  3815 => std_logic_vector'(x"00000000"),
  3816 => std_logic_vector'(x"00000000"),
  3817 => std_logic_vector'(x"00000000"),
  3818 => std_logic_vector'(x"00000000"),
  3819 => std_logic_vector'(x"00000000"),
  3820 => std_logic_vector'(x"00000000"),
  3821 => std_logic_vector'(x"00000000"),
  3822 => std_logic_vector'(x"00000000"),
  3823 => std_logic_vector'(x"00000000"),
  3824 => std_logic_vector'(x"00000000"),
  3825 => std_logic_vector'(x"00000000"),
  3826 => std_logic_vector'(x"00000000"),
  3827 => std_logic_vector'(x"00000000"),
  3828 => std_logic_vector'(x"00000000"),
  3829 => std_logic_vector'(x"00000000"),
  3830 => std_logic_vector'(x"00000000"),
  3831 => std_logic_vector'(x"00000000"),
  3832 => std_logic_vector'(x"00000000"),
  3833 => std_logic_vector'(x"00000000"),
  3834 => std_logic_vector'(x"00000000"),
  3835 => std_logic_vector'(x"00000000"),
  3836 => std_logic_vector'(x"00000000"),
  3837 => std_logic_vector'(x"00000000"),
  3838 => std_logic_vector'(x"00000000"),
  3839 => std_logic_vector'(x"00000000"),
  3840 => std_logic_vector'(x"00000000"),
  3841 => std_logic_vector'(x"00000000"),
  3842 => std_logic_vector'(x"00000000"),
  3843 => std_logic_vector'(x"00000000"),
  3844 => std_logic_vector'(x"00000000"),
  3845 => std_logic_vector'(x"00000000"),
  3846 => std_logic_vector'(x"00000000"),
  3847 => std_logic_vector'(x"00000000"),
  3848 => std_logic_vector'(x"00000000"),
  3849 => std_logic_vector'(x"00000000"),
  3850 => std_logic_vector'(x"00000000"),
  3851 => std_logic_vector'(x"00000000"),
  3852 => std_logic_vector'(x"00000000"),
  3853 => std_logic_vector'(x"00000000"),
  3854 => std_logic_vector'(x"00000000"),
  3855 => std_logic_vector'(x"00000000"),
  3856 => std_logic_vector'(x"00000000"),
  3857 => std_logic_vector'(x"00000000"),
  3858 => std_logic_vector'(x"00000000"),
  3859 => std_logic_vector'(x"00000000"),
  3860 => std_logic_vector'(x"00000000"),
  3861 => std_logic_vector'(x"00000000"),
  3862 => std_logic_vector'(x"00000000"),
  3863 => std_logic_vector'(x"00000000"),
  3864 => std_logic_vector'(x"00000000"),
  3865 => std_logic_vector'(x"00000000"),
  3866 => std_logic_vector'(x"00000000"),
  3867 => std_logic_vector'(x"00000000"),
  3868 => std_logic_vector'(x"00000000"),
  3869 => std_logic_vector'(x"00000000"),
  3870 => std_logic_vector'(x"00000000"),
  3871 => std_logic_vector'(x"00000000"),
  3872 => std_logic_vector'(x"00000000"),
  3873 => std_logic_vector'(x"00000000"),
  3874 => std_logic_vector'(x"00000000"),
  3875 => std_logic_vector'(x"00000000"),
  3876 => std_logic_vector'(x"00000000"),
  3877 => std_logic_vector'(x"00000000"),
  3878 => std_logic_vector'(x"00000000"),
  3879 => std_logic_vector'(x"00000000"),
  3880 => std_logic_vector'(x"00000000"),
  3881 => std_logic_vector'(x"00000000"),
  3882 => std_logic_vector'(x"00000000"),
  3883 => std_logic_vector'(x"00000000"),
  3884 => std_logic_vector'(x"00000000"),
  3885 => std_logic_vector'(x"00000000"),
  3886 => std_logic_vector'(x"00000000"),
  3887 => std_logic_vector'(x"00000000"),
  3888 => std_logic_vector'(x"00000000"),
  3889 => std_logic_vector'(x"00000000"),
  3890 => std_logic_vector'(x"00000000"),
  3891 => std_logic_vector'(x"00000000"),
  3892 => std_logic_vector'(x"00000000"),
  3893 => std_logic_vector'(x"00000000"),
  3894 => std_logic_vector'(x"00000000"),
  3895 => std_logic_vector'(x"00000000"),
  3896 => std_logic_vector'(x"00000000"),
  3897 => std_logic_vector'(x"00000000"),
  3898 => std_logic_vector'(x"00000000"),
  3899 => std_logic_vector'(x"00000000"),
  3900 => std_logic_vector'(x"00000000"),
  3901 => std_logic_vector'(x"00000000"),
  3902 => std_logic_vector'(x"00000000"),
  3903 => std_logic_vector'(x"00000000"),
  3904 => std_logic_vector'(x"00000000"),
  3905 => std_logic_vector'(x"00000000"),
  3906 => std_logic_vector'(x"00000000"),
  3907 => std_logic_vector'(x"00000000"),
  3908 => std_logic_vector'(x"00000000"),
  3909 => std_logic_vector'(x"00000000"),
  3910 => std_logic_vector'(x"00000000"),
  3911 => std_logic_vector'(x"00000000"),
  3912 => std_logic_vector'(x"00000000"),
  3913 => std_logic_vector'(x"00000000"),
  3914 => std_logic_vector'(x"00000000"),
  3915 => std_logic_vector'(x"00000000"),
  3916 => std_logic_vector'(x"00000000"),
  3917 => std_logic_vector'(x"00000000"),
  3918 => std_logic_vector'(x"00000000"),
  3919 => std_logic_vector'(x"00000000"),
  3920 => std_logic_vector'(x"00000000"),
  3921 => std_logic_vector'(x"00000000"),
  3922 => std_logic_vector'(x"00000000"),
  3923 => std_logic_vector'(x"00000000"),
  3924 => std_logic_vector'(x"00000000"),
  3925 => std_logic_vector'(x"00000000"),
  3926 => std_logic_vector'(x"00000000"),
  3927 => std_logic_vector'(x"00000000"),
  3928 => std_logic_vector'(x"00000000"),
  3929 => std_logic_vector'(x"00000000"),
  3930 => std_logic_vector'(x"00000000"),
  3931 => std_logic_vector'(x"00000000"),
  3932 => std_logic_vector'(x"00000000"),
  3933 => std_logic_vector'(x"00000000"),
  3934 => std_logic_vector'(x"00000000"),
  3935 => std_logic_vector'(x"00000000"),
  3936 => std_logic_vector'(x"00000000"),
  3937 => std_logic_vector'(x"00000000"),
  3938 => std_logic_vector'(x"00000000"),
  3939 => std_logic_vector'(x"00000000"),
  3940 => std_logic_vector'(x"00000000"),
  3941 => std_logic_vector'(x"00000000"),
  3942 => std_logic_vector'(x"00000000"),
  3943 => std_logic_vector'(x"00000000"),
  3944 => std_logic_vector'(x"00000000"),
  3945 => std_logic_vector'(x"00000000"),
  3946 => std_logic_vector'(x"00000000"),
  3947 => std_logic_vector'(x"00000000"),
  3948 => std_logic_vector'(x"00000000"),
  3949 => std_logic_vector'(x"00000000"),
  3950 => std_logic_vector'(x"00000000"),
  3951 => std_logic_vector'(x"00000000"),
  3952 => std_logic_vector'(x"00000000"),
  3953 => std_logic_vector'(x"00000000"),
  3954 => std_logic_vector'(x"00000000"),
  3955 => std_logic_vector'(x"00000000"),
  3956 => std_logic_vector'(x"00000000"),
  3957 => std_logic_vector'(x"00000000"),
  3958 => std_logic_vector'(x"00000000"),
  3959 => std_logic_vector'(x"00000000"),
  3960 => std_logic_vector'(x"00000000"),
  3961 => std_logic_vector'(x"00000000"),
  3962 => std_logic_vector'(x"00000000"),
  3963 => std_logic_vector'(x"00000000"),
  3964 => std_logic_vector'(x"00000000"),
  3965 => std_logic_vector'(x"00000000"),
  3966 => std_logic_vector'(x"00000000"),
  3967 => std_logic_vector'(x"00000000"),
  3968 => std_logic_vector'(x"00000000"),
  3969 => std_logic_vector'(x"00000000"),
  3970 => std_logic_vector'(x"00000000"),
  3971 => std_logic_vector'(x"00000000"),
  3972 => std_logic_vector'(x"00000000"),
  3973 => std_logic_vector'(x"00000000"),
  3974 => std_logic_vector'(x"00000000"),
  3975 => std_logic_vector'(x"00000000"),
  3976 => std_logic_vector'(x"00000000"),
  3977 => std_logic_vector'(x"00000000"),
  3978 => std_logic_vector'(x"00000000"),
  3979 => std_logic_vector'(x"00000000"),
  3980 => std_logic_vector'(x"00000000"),
  3981 => std_logic_vector'(x"00000000"),
  3982 => std_logic_vector'(x"00000000"),
  3983 => std_logic_vector'(x"00000000"),
  3984 => std_logic_vector'(x"00000000"),
  3985 => std_logic_vector'(x"00000000"),
  3986 => std_logic_vector'(x"00000000"),
  3987 => std_logic_vector'(x"00000000"),
  3988 => std_logic_vector'(x"00000000"),
  3989 => std_logic_vector'(x"00000000"),
  3990 => std_logic_vector'(x"00000000"),
  3991 => std_logic_vector'(x"00000000"),
  3992 => std_logic_vector'(x"00000000"),
  3993 => std_logic_vector'(x"00000000"),
  3994 => std_logic_vector'(x"00000000"),
  3995 => std_logic_vector'(x"00000000"),
  3996 => std_logic_vector'(x"00000000"),
  3997 => std_logic_vector'(x"00000000"),
  3998 => std_logic_vector'(x"00000000"),
  3999 => std_logic_vector'(x"00000000"),
  4000 => std_logic_vector'(x"00000000"),
  4001 => std_logic_vector'(x"00000000"),
  4002 => std_logic_vector'(x"00000000"),
  4003 => std_logic_vector'(x"00000000"),
  4004 => std_logic_vector'(x"00000000"),
  4005 => std_logic_vector'(x"00000000"),
  4006 => std_logic_vector'(x"00000000"),
  4007 => std_logic_vector'(x"00000000"),
  4008 => std_logic_vector'(x"00000000"),
  4009 => std_logic_vector'(x"00000000"),
  4010 => std_logic_vector'(x"00000000"),
  4011 => std_logic_vector'(x"00000000"),
  4012 => std_logic_vector'(x"00000000"),
  4013 => std_logic_vector'(x"00000000"),
  4014 => std_logic_vector'(x"00000000"),
  4015 => std_logic_vector'(x"00000000"),
  4016 => std_logic_vector'(x"00000000"),
  4017 => std_logic_vector'(x"00000000"),
  4018 => std_logic_vector'(x"00000000"),
  4019 => std_logic_vector'(x"00000000"),
  4020 => std_logic_vector'(x"00000000"),
  4021 => std_logic_vector'(x"00000000"),
  4022 => std_logic_vector'(x"00000000"),
  4023 => std_logic_vector'(x"00000000"),
  4024 => std_logic_vector'(x"00000000"),
  4025 => std_logic_vector'(x"00000000"),
  4026 => std_logic_vector'(x"00000000"),
  4027 => std_logic_vector'(x"00000000"),
  4028 => std_logic_vector'(x"00000000"),
  4029 => std_logic_vector'(x"00000000"),
  4030 => std_logic_vector'(x"00000000"),
  4031 => std_logic_vector'(x"00000000"),
  4032 => std_logic_vector'(x"00000000"),
  4033 => std_logic_vector'(x"00000000"),
  4034 => std_logic_vector'(x"00000000"),
  4035 => std_logic_vector'(x"00000000"),
  4036 => std_logic_vector'(x"00000000"),
  4037 => std_logic_vector'(x"00000000"),
  4038 => std_logic_vector'(x"00000000"),
  4039 => std_logic_vector'(x"00000000"),
  4040 => std_logic_vector'(x"00000000"),
  4041 => std_logic_vector'(x"00000000"),
  4042 => std_logic_vector'(x"00000000"),
  4043 => std_logic_vector'(x"00000000"),
  4044 => std_logic_vector'(x"00000000"),
  4045 => std_logic_vector'(x"00000000"),
  4046 => std_logic_vector'(x"00000000"),
  4047 => std_logic_vector'(x"00000000"),
  4048 => std_logic_vector'(x"00000000"),
  4049 => std_logic_vector'(x"00000000"),
  4050 => std_logic_vector'(x"00000000"),
  4051 => std_logic_vector'(x"00000000"),
  4052 => std_logic_vector'(x"00000000"),
  4053 => std_logic_vector'(x"00000000"),
  4054 => std_logic_vector'(x"00000000"),
  4055 => std_logic_vector'(x"00000000"),
  4056 => std_logic_vector'(x"00000000"),
  4057 => std_logic_vector'(x"00000000"),
  4058 => std_logic_vector'(x"00000000"),
  4059 => std_logic_vector'(x"00000000"),
  4060 => std_logic_vector'(x"00000000"),
  4061 => std_logic_vector'(x"00000000"),
  4062 => std_logic_vector'(x"00000000"),
  4063 => std_logic_vector'(x"00000000"),
  4064 => std_logic_vector'(x"00000000"),
  4065 => std_logic_vector'(x"00000000"),
  4066 => std_logic_vector'(x"00000000"),
  4067 => std_logic_vector'(x"00000000"),
  4068 => std_logic_vector'(x"00000000"),
  4069 => std_logic_vector'(x"00000000"),
  4070 => std_logic_vector'(x"00000000"),
  4071 => std_logic_vector'(x"00000000"),
  4072 => std_logic_vector'(x"00000000"),
  4073 => std_logic_vector'(x"00000000"),
  4074 => std_logic_vector'(x"00000000"),
  4075 => std_logic_vector'(x"00000000"),
  4076 => std_logic_vector'(x"00000000"),
  4077 => std_logic_vector'(x"00000000"),
  4078 => std_logic_vector'(x"00000000"),
  4079 => std_logic_vector'(x"00000000"),
  4080 => std_logic_vector'(x"00000000"),
  4081 => std_logic_vector'(x"00000000"),
  4082 => std_logic_vector'(x"00000000"),
  4083 => std_logic_vector'(x"00000000"),
  4084 => std_logic_vector'(x"00000000"),
  4085 => std_logic_vector'(x"00000000"),
  4086 => std_logic_vector'(x"00000000"),
  4087 => std_logic_vector'(x"00000000"),
  4088 => std_logic_vector'(x"00000000"),
  4089 => std_logic_vector'(x"00000000"),
  4090 => std_logic_vector'(x"00000000"),
  4091 => std_logic_vector'(x"00000000"),
  4092 => std_logic_vector'(x"00000000"),
  4093 => std_logic_vector'(x"00000000"),
  4094 => std_logic_vector'(x"00000000"),
  4095 => std_logic_vector'(x"00000000"),
  4096 => std_logic_vector'(x"31020000"),
  4097 => std_logic_vector'(x"0004002b"),
  4098 => std_logic_vector'(x"31024000"),
  4099 => std_logic_vector'(x"0008002d"),
  4100 => std_logic_vector'(x"30024008"),
  4101 => std_logic_vector'(x"000e003d"),
  4102 => std_logic_vector'(x"63054010"),
  4103 => std_logic_vector'(x"2b6c6c65"),
  4104 => std_logic_vector'(x"40180012"),
  4105 => std_logic_vector'(x"6c656305"),
  4106 => std_logic_vector'(x"0016736c"),
  4107 => std_logic_vector'(x"3c024022"),
  4108 => std_logic_vector'(x"001a003e"),
  4109 => std_logic_vector'(x"3e01402c"),
  4110 => std_logic_vector'(x"4034001e"),
  4111 => std_logic_vector'(x"003c3002"),
  4112 => std_logic_vector'(x"403a0022"),
  4113 => std_logic_vector'(x"003e3002"),
  4114 => std_logic_vector'(x"40420026"),
  4115 => std_logic_vector'(x"3e3c3003"),
  4116 => std_logic_vector'(x"404a002a"),
  4117 => std_logic_vector'(x"003e7502"),
  4118 => std_logic_vector'(x"4052002e"),
  4119 => std_logic_vector'(x"79656b04"),
  4120 => std_logic_vector'(x"003a003f"),
  4121 => std_logic_vector'(x"6b03405a"),
  4122 => std_logic_vector'(x"00467965"),
  4123 => std_logic_vector'(x"65044064"),
  4124 => std_logic_vector'(x"0074696d"),
  4125 => std_logic_vector'(x"406c0050"),
  4126 => std_logic_vector'(x"00726302"),
  4127 => std_logic_vector'(x"4076005c"),
  4128 => std_logic_vector'(x"61707305"),
  4129 => std_logic_vector'(x"00646563"),
  4130 => std_logic_vector'(x"6202407e"),
  4131 => std_logic_vector'(x"0068006c"),
  4132 => std_logic_vector'(x"2e024088"),
  4133 => std_logic_vector'(x"009a0078"),
  4134 => std_logic_vector'(x"66054090"),
  4135 => std_logic_vector'(x"65736c61"),
  4136 => std_logic_vector'(x"4098009e"),
  4137 => std_logic_vector'(x"75727404"),
  4138 => std_logic_vector'(x"00a20065"),
  4139 => std_logic_vector'(x"720340a2"),
  4140 => std_logic_vector'(x"00a6746f"),
  4141 => std_logic_vector'(x"2d0440ac"),
  4142 => std_logic_vector'(x"00746f72"),
  4143 => std_logic_vector'(x"40b400ae"),
  4144 => std_logic_vector'(x"63757404"),
  4145 => std_logic_vector'(x"00b8006b"),
  4146 => std_logic_vector'(x"320540be"),
  4147 => std_logic_vector'(x"706f7264"),
  4148 => std_logic_vector'(x"40c800bc"),
  4149 => std_logic_vector'(x"75643f04"),
  4150 => std_logic_vector'(x"00c00070"),
  4151 => std_logic_vector'(x"320440d2"),
  4152 => std_logic_vector'(x"00707564"),
  4153 => std_logic_vector'(x"40dc00c8"),
  4154 => std_logic_vector'(x"00212b02"),
  4155 => std_logic_vector'(x"40e600cc"),
  4156 => std_logic_vector'(x"77733205"),
  4157 => std_logic_vector'(x"00da7061"),
  4158 => std_logic_vector'(x"320540ee"),
  4159 => std_logic_vector'(x"7265766f"),
  4160 => std_logic_vector'(x"40f800e4"),
  4161 => std_logic_vector'(x"6e696d03"),
  4162 => std_logic_vector'(x"410200f0"),
  4163 => std_logic_vector'(x"78616d03"),
  4164 => std_logic_vector'(x"410a00fc"),
  4165 => std_logic_vector'(x"00406302"),
  4166 => std_logic_vector'(x"41120108"),
  4167 => std_logic_vector'(x"40777503"),
  4168 => std_logic_vector'(x"411a0126"),
  4169 => std_logic_vector'(x"00407702"),
  4170 => std_logic_vector'(x"41220136"),
  4171 => std_logic_vector'(x"00217702"),
  4172 => std_logic_vector'(x"412a0156"),
  4173 => std_logic_vector'(x"00216302"),
  4174 => std_logic_vector'(x"41320188"),
  4175 => std_logic_vector'(x"756f6305"),
  4176 => std_logic_vector'(x"01b2746e"),
  4177 => std_logic_vector'(x"6206413a"),
  4178 => std_logic_vector'(x"646e756f"),
  4179 => std_logic_vector'(x"01ba0073"),
  4180 => std_logic_vector'(x"74044144"),
  4181 => std_logic_vector'(x"00657079"),
  4182 => std_logic_vector'(x"000001c0"),
  4183 => std_logic_vector'(x"646c6f63"),
  4184 => std_logic_vector'(x"00000010"),
  4185 => std_logic_vector'(x"00005606"),
  4186 => std_logic_vector'(x"000023ea"),
  4187 => std_logic_vector'(x"00005618"),
  4188 => std_logic_vector'(x"00005606"),
  4189 => std_logic_vector'(x"000023dc"),
  4190 => std_logic_vector'(x"000023dc"),
  4191 => std_logic_vector'(x"0000002a"),
  4192 => std_logic_vector'(x"000041a0"),
  4193 => std_logic_vector'(x"00000000"),
  4194 => std_logic_vector'(x"00000009"),
  4195 => std_logic_vector'(x"00000000"),
  4196 => std_logic_vector'(x"00000029"),
  4197 => std_logic_vector'(x"00000000"),
  4198 => std_logic_vector'(x"00000000"),
  4199 => std_logic_vector'(x"00000001"),
  4200 => std_logic_vector'(x"35343332"),
  4201 => std_logic_vector'(x"406f6920"),
  4202 => std_logic_vector'(x"44205c20"),
  4203 => std_logic_vector'(x"20706d75"),
  4204 => std_logic_vector'(x"20656874"),
  4205 => std_logic_vector'(x"6f6d656d"),
  4206 => std_logic_vector'(x"74207972"),
  4207 => std_logic_vector'(x"656d206f"),
  4208 => std_logic_vector'(x"75645f6d"),
  4209 => std_logic_vector'(x"682e706d"),
  4210 => std_logic_vector'(x"74207865"),
  4211 => std_logic_vector'(x"62747365"),
  4212 => std_logic_vector'(x"68636e65"),
  4213 => std_logic_vector'(x"74697720"),
  4214 => std_logic_vector'(x"656d2068"),
  4215 => std_logic_vector'(x"79726f6d"),
  4216 => std_logic_vector'(x"6d756420"),
  4217 => std_logic_vector'(x"66207370"),
  4218 => std_logic_vector'(x"206d6f72"),
  4219 => std_logic_vector'(x"6e616863"),
  4220 => std_logic_vector'(x"206c656e"),
  4221 => std_logic_vector'(x"3c3c3130"),
  4222 => std_logic_vector'(x"69293831"),
  4223 => std_logic_vector'(x"6d206874"),
  4224 => std_logic_vector'(x"69746c75"),
  4225 => std_logic_vector'(x"20656c70"),
  4226 => std_logic_vector'(x"74697865"),
  4227 => std_logic_vector'(x"696f7020"),
  4228 => std_logic_vector'(x"6c73746e"),
  4229 => std_logic_vector'(x"77614220"),
  4230 => std_logic_vector'(x"00002e64"),
  4231 => std_logic_vector'(x"00000000"),
  4232 => std_logic_vector'(x"64024150"),
  4233 => std_logic_vector'(x"01d20070"),
  4234 => std_logic_vector'(x"63024220"),
  4235 => std_logic_vector'(x"01d60070"),
  4236 => std_logic_vector'(x"73054228"),
  4237 => std_logic_vector'(x"65746174"),
  4238 => std_logic_vector'(x"423001da"),
  4239 => std_logic_vector'(x"73616204"),
  4240 => std_logic_vector'(x"01de0065"),
  4241 => std_logic_vector'(x"3e03423a"),
  4242 => std_logic_vector'(x"01e26e69"),
  4243 => std_logic_vector'(x"66054244"),
  4244 => std_logic_vector'(x"6874726f"),
  4245 => std_logic_vector'(x"424c01e6"),
  4246 => std_logic_vector'(x"68747403"),
  4247 => std_logic_vector'(x"425601ea"),
  4248 => std_logic_vector'(x"726f7705"),
  4249 => std_logic_vector'(x"01f67364"),
  4250 => std_logic_vector'(x"6e06425e"),
  4251 => std_logic_vector'(x"74616765"),
  4252 => std_logic_vector'(x"02100065"),
  4253 => std_logic_vector'(x"2d014268"),
  4254 => std_logic_vector'(x"42740214"),
  4255 => std_logic_vector'(x"73626103"),
  4256 => std_logic_vector'(x"427a0218"),
  4257 => std_logic_vector'(x"002a3202"),
  4258 => std_logic_vector'(x"42820222"),
  4259 => std_logic_vector'(x"002f3202"),
  4260 => std_logic_vector'(x"428a0226"),
  4261 => std_logic_vector'(x"72656804"),
  4262 => std_logic_vector'(x"023c0065"),
  4263 => std_logic_vector'(x"64054292"),
  4264 => std_logic_vector'(x"68747065"),
  4265 => std_logic_vector'(x"429c0242"),
  4266 => std_logic_vector'(x"74732f07"),
  4267 => std_logic_vector'(x"676e6972"),
  4268 => std_logic_vector'(x"42a60248"),
  4269 => std_logic_vector'(x"696c6107"),
  4270 => std_logic_vector'(x"64656e67"),
  4271 => std_logic_vector'(x"42b20256"),
  4272 => std_logic_vector'(x"002b6402"),
  4273 => std_logic_vector'(x"42be0260"),
  4274 => std_logic_vector'(x"656e6407"),
  4275 => std_logic_vector'(x"65746167"),
  4276 => std_logic_vector'(x"42c6027c"),
  4277 => std_logic_vector'(x"62616404"),
  4278 => std_logic_vector'(x"028a0073"),
  4279 => std_logic_vector'(x"730342d2"),
  4280 => std_logic_vector'(x"0294643e"),
  4281 => std_logic_vector'(x"320242dc"),
  4282 => std_logic_vector'(x"02980040"),
  4283 => std_logic_vector'(x"320242e4"),
  4284 => std_logic_vector'(x"02a60021"),
  4285 => std_logic_vector'(x"320442ec"),
  4286 => std_logic_vector'(x"00746f72"),
  4287 => std_logic_vector'(x"42f402b2"),
  4288 => std_logic_vector'(x"733e6403"),
  4289 => std_logic_vector'(x"42fe02be"),
  4290 => std_logic_vector'(x"003d6402"),
  4291 => std_logic_vector'(x"430602c0"),
  4292 => std_logic_vector'(x"003c6402"),
  4293 => std_logic_vector'(x"430e02ce"),
  4294 => std_logic_vector'(x"3c756403"),
  4295 => std_logic_vector'(x"431602e4"),
  4296 => std_logic_vector'(x"002d6402"),
  4297 => std_logic_vector'(x"431e02fa"),
  4298 => std_logic_vector'(x"3c306403"),
  4299 => std_logic_vector'(x"432602fe"),
  4300 => std_logic_vector'(x"3d306403"),
  4301 => std_logic_vector'(x"432e0302"),
  4302 => std_logic_vector'(x"2a326403"),
  4303 => std_logic_vector'(x"43360306"),
  4304 => std_logic_vector'(x"2f326403"),
  4305 => std_logic_vector'(x"0000030a"),
  4306 => std_logic_vector'(x"00000010"),
  4307 => std_logic_vector'(x"7503433e"),
  4308 => std_logic_vector'(x"03542a6d"),
  4309 => std_logic_vector'(x"2a01434c"),
  4310 => std_logic_vector'(x"4354038a"),
  4311 => std_logic_vector'(x"2f6d7506"),
  4312 => std_logic_vector'(x"00646f6d"),
  4313 => std_logic_vector'(x"435a03ca"),
  4314 => std_logic_vector'(x"63636106"),
  4315 => std_logic_vector'(x"00747065"),
  4316 => std_logic_vector'(x"436603fc"),
  4317 => std_logic_vector'(x"6c616308"),
  4318 => std_logic_vector'(x"656e6769"),
  4319 => std_logic_vector'(x"04ea0064"),
  4320 => std_logic_vector'(x"63064372"),
  4321 => std_logic_vector'(x"67696c61"),
  4322 => std_logic_vector'(x"04fe006e"),
  4323 => std_logic_vector'(x"73054380"),
  4324 => std_logic_vector'(x"646e6966"),
  4325 => std_logic_vector'(x"438c0516"),
  4326 => std_logic_vector'(x"756e3e07"),
  4327 => std_logic_vector'(x"7265626d"),
  4328 => std_logic_vector'(x"4396056a"),
  4329 => std_logic_vector'(x"6c696604"),
  4330 => std_logic_vector'(x"0598006c"),
  4331 => std_logic_vector'(x"630543a2"),
  4332 => std_logic_vector'(x"65766f6d"),
  4333 => std_logic_vector'(x"43ac05b0"),
  4334 => std_logic_vector'(x"6f6d6306"),
  4335 => std_logic_vector'(x"003e6576"),
  4336 => std_logic_vector'(x"43b605d0"),
  4337 => std_logic_vector'(x"65786507"),
  4338 => std_logic_vector'(x"65747563"),
  4339 => std_logic_vector'(x"43c205f0"),
  4340 => std_logic_vector'(x"756f7306"),
  4341 => std_logic_vector'(x"00656372"),
  4342 => std_logic_vector'(x"43ce05f4"),
  4343 => std_logic_vector'(x"756f7309"),
  4344 => std_logic_vector'(x"2d656372"),
  4345 => std_logic_vector'(x"05fc6469"),
  4346 => std_logic_vector'(x"700a43da"),
  4347 => std_logic_vector'(x"65737261"),
  4348 => std_logic_vector'(x"6d616e2d"),
  4349 => std_logic_vector'(x"06220065"),
  4350 => std_logic_vector'(x"700543e8"),
  4351 => std_logic_vector'(x"65737261"),
  4352 => std_logic_vector'(x"43f8065c"),
  4353 => std_logic_vector'(x"6c6c6105"),
  4354 => std_logic_vector'(x"0690746f"),
  4355 => std_logic_vector'(x"2c014402"),
  4356 => std_logic_vector'(x"440c0694"),
  4357 => std_logic_vector'(x"002c7702"),
  4358 => std_logic_vector'(x"4412069e"),
  4359 => std_logic_vector'(x"002c6302"),
  4360 => std_logic_vector'(x"441a06a6"),
  4361 => std_logic_vector'(x"002c7302"),
  4362 => std_logic_vector'(x"442206da"),
  4363 => std_logic_vector'(x"6d6d6909"),
  4364 => std_logic_vector'(x"61696465"),
  4365 => std_logic_vector'(x"071a6574"),
  4366 => std_logic_vector'(x"5d01442a"),
  4367 => std_logic_vector'(x"4439072c"),
  4368 => std_logic_vector'(x"07345b01"),
  4369 => std_logic_vector'(x"3a01443e"),
  4370 => std_logic_vector'(x"4444073c"),
  4371 => std_logic_vector'(x"6f6e3a07"),
  4372 => std_logic_vector'(x"656d616e"),
  4373 => std_logic_vector'(x"444b0740"),
  4374 => std_logic_vector'(x"69786504"),
  4375 => std_logic_vector'(x"07a80074"),
  4376 => std_logic_vector'(x"3b014457"),
  4377 => std_logic_vector'(x"446107d8"),
  4378 => std_logic_vector'(x"00666902"),
  4379 => std_logic_vector'(x"446707de"),
  4380 => std_logic_vector'(x"65686105"),
  4381 => std_logic_vector'(x"07e86461"),
  4382 => std_logic_vector'(x"7404446f"),
  4383 => std_logic_vector'(x"006e6568"),
  4384 => std_logic_vector'(x"447907f2"),
  4385 => std_logic_vector'(x"67656205"),
  4386 => std_logic_vector'(x"08066e69"),
  4387 => std_logic_vector'(x"61054483"),
  4388 => std_logic_vector'(x"6e696167"),
  4389 => std_logic_vector'(x"448d080e"),
  4390 => std_logic_vector'(x"746e7505"),
  4391 => std_logic_vector'(x"08106c69"),
  4392 => std_logic_vector'(x"63084496"),
  4393 => std_logic_vector'(x"69706d6f"),
  4394 => std_logic_vector'(x"002c656c"),
  4395 => std_logic_vector'(x"44a00846"),
  4396 => std_logic_vector'(x"656f6405"),
  4397 => std_logic_vector'(x"08763e73"),
  4398 => std_logic_vector'(x"720744af"),
  4399 => std_logic_vector'(x"72756365"),
  4400 => std_logic_vector'(x"08886573"),
  4401 => std_logic_vector'(x"640244b9"),
  4402 => std_logic_vector'(x"08ca006f"),
  4403 => std_logic_vector'(x"6c0444c5"),
  4404 => std_logic_vector'(x"00706f6f"),
  4405 => std_logic_vector'(x"44cd090e"),
  4406 => std_logic_vector'(x"6f6c2b05"),
  4407 => std_logic_vector'(x"093e706f"),
  4408 => std_logic_vector'(x"6c0544d7"),
  4409 => std_logic_vector'(x"65766165"),
  4410 => std_logic_vector'(x"44e1094a"),
  4411 => std_logic_vector'(x"6f643f03"),
  4412 => std_logic_vector'(x"44ea0962"),
  4413 => std_logic_vector'(x"09946901"),
  4414 => std_logic_vector'(x"6a0144f2"),
  4415 => std_logic_vector'(x"44f909a6"),
  4416 => std_logic_vector'(x"6c6e7506"),
  4417 => std_logic_vector'(x"00706f6f"),
  4418 => std_logic_vector'(x"44fe09c0"),
  4419 => std_logic_vector'(x"63656407"),
  4420 => std_logic_vector'(x"6c616d69"),
  4421 => std_logic_vector'(x"450a09c8"),
  4422 => std_logic_vector'(x"09d02101"),
  4423 => std_logic_vector'(x"2b014516"),
  4424 => std_logic_vector'(x"451c09d4"),
  4425 => std_logic_vector'(x"726f7803"),
  4426 => std_logic_vector'(x"452209d6"),
  4427 => std_logic_vector'(x"646e6103"),
  4428 => std_logic_vector'(x"452a09d8"),
  4429 => std_logic_vector'(x"00726f02"),
  4430 => std_logic_vector'(x"453209da"),
  4431 => std_logic_vector'(x"766e6906"),
  4432 => std_logic_vector'(x"00747265"),
  4433 => std_logic_vector'(x"453a09dc"),
  4434 => std_logic_vector'(x"09de3d01"),
  4435 => std_logic_vector'(x"3c014546"),
  4436 => std_logic_vector'(x"454c09e0"),
  4437 => std_logic_vector'(x"003c7502"),
  4438 => std_logic_vector'(x"455209e2"),
  4439 => std_logic_vector'(x"61777304"),
  4440 => std_logic_vector'(x"09e40070"),
  4441 => std_logic_vector'(x"6403455a"),
  4442 => std_logic_vector'(x"09e67075"),
  4443 => std_logic_vector'(x"64044564"),
  4444 => std_logic_vector'(x"00706f72"),
  4445 => std_logic_vector'(x"456c09e8"),
  4446 => std_logic_vector'(x"65766f04"),
  4447 => std_logic_vector'(x"09ea0072"),
  4448 => std_logic_vector'(x"6e034576"),
  4449 => std_logic_vector'(x"09ec7069"),
  4450 => std_logic_vector'(x"40014580"),
  4451 => std_logic_vector'(x"458809ee"),
  4452 => std_logic_vector'(x"216f6903"),
  4453 => std_logic_vector'(x"458e09f2"),
  4454 => std_logic_vector'(x"406f6903"),
  4455 => std_logic_vector'(x"459609f6"),
  4456 => std_logic_vector'(x"68737206"),
  4457 => std_logic_vector'(x"00746669"),
  4458 => std_logic_vector'(x"459e09fa"),
  4459 => std_logic_vector'(x"68736c06"),
  4460 => std_logic_vector'(x"00746669"),
  4461 => std_logic_vector'(x"45ab09fc"),
  4462 => std_logic_vector'(x"00723e02"),
  4463 => std_logic_vector'(x"45b709fe"),
  4464 => std_logic_vector'(x"003e7202"),
  4465 => std_logic_vector'(x"45bf0a04"),
  4466 => std_logic_vector'(x"00407202"),
  4467 => std_logic_vector'(x"45c60a0a"),
  4468 => std_logic_vector'(x"72687405"),
  4469 => std_logic_vector'(x"0a18776f"),
  4470 => std_logic_vector'(x"320845cf"),
  4471 => std_logic_vector'(x"6574696c"),
  4472 => std_logic_vector'(x"006c6172"),
  4473 => std_logic_vector'(x"45d90a44"),
  4474 => std_logic_vector'(x"74696c07"),
  4475 => std_logic_vector'(x"6c617265"),
  4476 => std_logic_vector'(x"45e70a48"),
  4477 => std_logic_vector'(x"736f7008"),
  4478 => std_logic_vector'(x"6e6f7074"),
  4479 => std_logic_vector'(x"0b460065"),
  4480 => std_logic_vector'(x"720645f2"),
  4481 => std_logic_vector'(x"6c696665"),
  4482 => std_logic_vector'(x"0b88006c"),
  4483 => std_logic_vector'(x"65084600"),
  4484 => std_logic_vector'(x"756c6176"),
  4485 => std_logic_vector'(x"00657461"),
  4486 => std_logic_vector'(x"460c0ba4"),
  4487 => std_logic_vector'(x"69757104"),
  4488 => std_logic_vector'(x"0be20074"),
  4489 => std_logic_vector'(x"0000461a"),
  4490 => std_logic_vector'(x"5c01461b"),
  4491 => std_logic_vector'(x"46280c0e"),
  4492 => std_logic_vector'(x"61686305"),
  4493 => std_logic_vector'(x"0c182b72"),
  4494 => std_logic_vector'(x"6305462e"),
  4495 => std_logic_vector'(x"73726168"),
  4496 => std_logic_vector'(x"46380c1c"),
  4497 => std_logic_vector'(x"6f626105"),
  4498 => std_logic_vector'(x"0c1e7472"),
  4499 => std_logic_vector'(x"27014642"),
  4500 => std_logic_vector'(x"464d0c26"),
  4501 => std_logic_vector'(x"5d275b03"),
  4502 => std_logic_vector'(x"46520c36"),
  4503 => std_logic_vector'(x"61686304"),
  4504 => std_logic_vector'(x"0c3c0072"),
  4505 => std_logic_vector'(x"5b06465b"),
  4506 => std_logic_vector'(x"72616863"),
  4507 => std_logic_vector'(x"0c44005d"),
  4508 => std_logic_vector'(x"28014665"),
  4509 => std_logic_vector'(x"46710c4a"),
  4510 => std_logic_vector'(x"736c6504"),
  4511 => std_logic_vector'(x"0c520065"),
  4512 => std_logic_vector'(x"77054677"),
  4513 => std_logic_vector'(x"656c6968"),
  4514 => std_logic_vector'(x"46810c5a"),
  4515 => std_logic_vector'(x"70657206"),
  4516 => std_logic_vector'(x"00746165"),
  4517 => std_logic_vector'(x"468a0c60"),
  4518 => std_logic_vector'(x"696c6105"),
  4519 => std_logic_vector'(x"0c666e67"),
  4520 => std_logic_vector'(x"32034696"),
  4521 => std_logic_vector'(x"0c70723e"),
  4522 => std_logic_vector'(x"320346a1"),
  4523 => std_logic_vector'(x"0c7e3e72"),
  4524 => std_logic_vector'(x"320346a8"),
  4525 => std_logic_vector'(x"0c884072"),
  4526 => std_logic_vector'(x"630646b0"),
  4527 => std_logic_vector'(x"74616572"),
  4528 => std_logic_vector'(x"0c9a0065"),
  4529 => std_logic_vector'(x"3e0546b8"),
  4530 => std_logic_vector'(x"79646f62"),
  4531 => std_logic_vector'(x"46c40ca6"),
  4532 => std_logic_vector'(x"61763209"),
  4533 => std_logic_vector'(x"62616972"),
  4534 => std_logic_vector'(x"0cae656c"),
  4535 => std_logic_vector'(x"320946ce"),
  4536 => std_logic_vector'(x"736e6f63"),
  4537 => std_logic_vector'(x"746e6174"),
  4538 => std_logic_vector'(x"46dc0cb8"),
  4539 => std_logic_vector'(x"616d6404"),
  4540 => std_logic_vector'(x"0cc40078"),
  4541 => std_logic_vector'(x"640446ea"),
  4542 => std_logic_vector'(x"006e696d"),
  4543 => std_logic_vector'(x"46f40cd2"),
  4544 => std_logic_vector'(x"002b6d02"),
  4545 => std_logic_vector'(x"46fe0ce2"),
  4546 => std_logic_vector'(x"002a6d02"),
  4547 => std_logic_vector'(x"47060ce8"),
  4548 => std_logic_vector'(x"656e7407"),
  4549 => std_logic_vector'(x"65746167"),
  4550 => std_logic_vector'(x"470e0d00"),
  4551 => std_logic_vector'(x"002a7402"),
  4552 => std_logic_vector'(x"471a0d18"),
  4553 => std_logic_vector'(x"002f7402"),
  4554 => std_logic_vector'(x"47220d42"),
  4555 => std_logic_vector'(x"2f2a6d03"),
  4556 => std_logic_vector'(x"472a0d6a"),
  4557 => std_logic_vector'(x"72617608"),
  4558 => std_logic_vector'(x"6c626169"),
  4559 => std_logic_vector'(x"0d740065"),
  4560 => std_logic_vector'(x"63084732"),
  4561 => std_logic_vector'(x"74736e6f"),
  4562 => std_logic_vector'(x"00746e61"),
  4563 => std_logic_vector'(x"47400d7c"),
  4564 => std_logic_vector'(x"6e677303"),
  4565 => std_logic_vector'(x"474e0d84"),
  4566 => std_logic_vector'(x"2f6d7306"),
  4567 => std_logic_vector'(x"006d6572"),
  4568 => std_logic_vector'(x"47560d8c"),
  4569 => std_logic_vector'(x"2f6d6606"),
  4570 => std_logic_vector'(x"00646f6d"),
  4571 => std_logic_vector'(x"47620dae"),
  4572 => std_logic_vector'(x"6d2f2a05"),
  4573 => std_logic_vector'(x"0dea646f"),
  4574 => std_logic_vector'(x"2a02476e"),
  4575 => std_logic_vector'(x"0df4002f"),
  4576 => std_logic_vector'(x"73064778"),
  4577 => std_logic_vector'(x"65636170"),
  4578 => std_logic_vector'(x"0dfa0073"),
  4579 => std_logic_vector'(x"42044780"),
  4580 => std_logic_vector'(x"00304655"),
  4581 => std_logic_vector'(x"00000e0a"),
  4582 => std_logic_vector'(x"00000000"),
  4583 => std_logic_vector'(x"00000000"),
  4584 => std_logic_vector'(x"00000000"),
  4585 => std_logic_vector'(x"00000000"),
  4586 => std_logic_vector'(x"00000000"),
  4587 => std_logic_vector'(x"00000000"),
  4588 => std_logic_vector'(x"00000000"),
  4589 => std_logic_vector'(x"00000000"),
  4590 => std_logic_vector'(x"00000000"),
  4591 => std_logic_vector'(x"00000000"),
  4592 => std_logic_vector'(x"00000000"),
  4593 => std_logic_vector'(x"00000000"),
  4594 => std_logic_vector'(x"00000000"),
  4595 => std_logic_vector'(x"00000000"),
  4596 => std_logic_vector'(x"00000000"),
  4597 => std_logic_vector'(x"00000000"),
  4598 => std_logic_vector'(x"478c0000"),
  4599 => std_logic_vector'(x"46554203"),
  4600 => std_logic_vector'(x"47da0e0e"),
  4601 => std_logic_vector'(x"646c6803"),
  4602 => std_logic_vector'(x"00000e12"),
  4603 => std_logic_vector'(x"00000000"),
  4604 => std_logic_vector'(x"3c0247e2"),
  4605 => std_logic_vector'(x"0e160023"),
  4606 => std_logic_vector'(x"680447f0"),
  4607 => std_logic_vector'(x"00646c6f"),
  4608 => std_logic_vector'(x"47f80e1e"),
  4609 => std_logic_vector'(x"67697304"),
  4610 => std_logic_vector'(x"0e2e006e"),
  4611 => std_logic_vector'(x"23014802"),
  4612 => std_logic_vector'(x"480c0e38"),
  4613 => std_logic_vector'(x"00732302"),
  4614 => std_logic_vector'(x"48120e60"),
  4615 => std_logic_vector'(x"003e2302"),
  4616 => std_logic_vector'(x"481a0e6a"),
  4617 => std_logic_vector'(x"722e6403"),
  4618 => std_logic_vector'(x"48220e78"),
  4619 => std_logic_vector'(x"002e6402"),
  4620 => std_logic_vector'(x"482a0e96"),
  4621 => std_logic_vector'(x"0e9e2e01"),
  4622 => std_logic_vector'(x"75024832"),
  4623 => std_logic_vector'(x"0ea4002e"),
  4624 => std_logic_vector'(x"2e024838"),
  4625 => std_logic_vector'(x"0eaa0072"),
  4626 => std_logic_vector'(x"75034840"),
  4627 => std_logic_vector'(x"0eb4722e"),
  4628 => std_logic_vector'(x"6d044848"),
  4629 => std_logic_vector'(x"0065766f"),
  4630 => std_logic_vector'(x"48500ebc"),
  4631 => std_logic_vector'(x"726f7704"),
  4632 => std_logic_vector'(x"0ed00064"),
  4633 => std_logic_vector'(x"2f04485a"),
  4634 => std_logic_vector'(x"00646f6d"),
  4635 => std_logic_vector'(x"48640f08"),
  4636 => std_logic_vector'(x"0f122f01"),
  4637 => std_logic_vector'(x"6d03486e"),
  4638 => std_logic_vector'(x"0f18646f"),
  4639 => std_logic_vector'(x"63024875"),
  4640 => std_logic_vector'(x"0f1e0022"),
  4641 => std_logic_vector'(x"7308487d"),
  4642 => std_logic_vector'(x"6574696c"),
  4643 => std_logic_vector'(x"006c6172"),
  4644 => std_logic_vector'(x"48840f2a"),
  4645 => std_logic_vector'(x"222e2804"),
  4646 => std_logic_vector'(x"0f360029"),
  4647 => std_logic_vector'(x"2e024893"),
  4648 => std_logic_vector'(x"0f3c0022"),
  4649 => std_logic_vector'(x"7506489c"),
  4650 => std_logic_vector'(x"6573756e"),
  4651 => std_logic_vector'(x"0f560064"),
  4652 => std_logic_vector'(x"700348a4"),
  4653 => std_logic_vector'(x"0f706461"),
  4654 => std_logic_vector'(x"720448b0"),
  4655 => std_logic_vector'(x"006c6c6f"),
  4656 => std_logic_vector'(x"48b80f76"),
  4657 => std_logic_vector'(x"63697004"),
  4658 => std_logic_vector'(x"0f88006b"),
  4659 => std_logic_vector'(x"650548c2"),
  4660 => std_logic_vector'(x"65736172"),
  4661 => std_logic_vector'(x"48cc0f9e"),
  4662 => std_logic_vector'(x"74697706"),
  4663 => std_logic_vector'(x"006e6968"),
  4664 => std_logic_vector'(x"48d70fa4"),
  4665 => std_logic_vector'(x"00282e02"),
  4666 => std_logic_vector'(x"48e20fb2"),
  4667 => std_logic_vector'(x"6e696604"),
  4668 => std_logic_vector'(x"0fba0064"),
  4669 => std_logic_vector'(x"5b0948eb"),
  4670 => std_logic_vector'(x"706d6f63"),
  4671 => std_logic_vector'(x"5d656c69"),
  4672 => std_logic_vector'(x"48f40fcc"),
  4673 => std_logic_vector'(x"0fd25f01"),
  4674 => std_logic_vector'(x"52312d64"),
  4675 => std_logic_vector'(x"5d545f44"),
  4676 => std_logic_vector'(x"00000000"),
  4677 => std_logic_vector'(x"00000000"),
  4678 => std_logic_vector'(x"00000000"),
  4679 => std_logic_vector'(x"00000000"),
  4680 => std_logic_vector'(x"00000000"),
  4681 => std_logic_vector'(x"00000000"),
  4682 => std_logic_vector'(x"00000000"),
  4683 => std_logic_vector'(x"00000000"),
  4684 => std_logic_vector'(x"00000000"),
  4685 => std_logic_vector'(x"00000000"),
  4686 => std_logic_vector'(x"00000000"),
  4687 => std_logic_vector'(x"00000000"),
  4688 => std_logic_vector'(x"00000000"),
  4689 => std_logic_vector'(x"00000000"),
  4690 => std_logic_vector'(x"00000000"),
  4691 => std_logic_vector'(x"00000000"),
  4692 => std_logic_vector'(x"00000000"),
  4693 => std_logic_vector'(x"00000000"),
  4694 => std_logic_vector'(x"73024903"),
  4695 => std_logic_vector'(x"0fd60022"),
  4696 => std_logic_vector'(x"63044959"),
  4697 => std_logic_vector'(x"00657361"),
  4698 => std_logic_vector'(x"49610ff2"),
  4699 => std_logic_vector'(x"00666f02"),
  4700 => std_logic_vector'(x"496b0ff6"),
  4701 => std_logic_vector'(x"646e6505"),
  4702 => std_logic_vector'(x"100a666f"),
  4703 => std_logic_vector'(x"65074973"),
  4704 => std_logic_vector'(x"6163646e"),
  4705 => std_logic_vector'(x"10126573"),
  4706 => std_logic_vector'(x"6803497c"),
  4707 => std_logic_vector'(x"10267865"),
  4708 => std_logic_vector'(x"730a4988"),
  4709 => std_logic_vector'(x"2d657661"),
  4710 => std_logic_vector'(x"75706e69"),
  4711 => std_logic_vector'(x"102e0074"),
  4712 => std_logic_vector'(x"720d4990"),
  4713 => std_logic_vector'(x"6f747365"),
  4714 => std_logic_vector'(x"692d6572"),
  4715 => std_logic_vector'(x"7475706e"),
  4716 => std_logic_vector'(x"49a01036"),
  4717 => std_logic_vector'(x"6e6f6307"),
  4718 => std_logic_vector'(x"74726576"),
  4719 => std_logic_vector'(x"49b21040"),
  4720 => std_logic_vector'(x"72616d06"),
  4721 => std_logic_vector'(x"0072656b"),
  4722 => std_logic_vector'(x"49be104a"),
  4723 => std_logic_vector'(x"74782e03"),
  4724 => std_logic_vector'(x"49ca107c"),
  4725 => std_logic_vector'(x"34706f03"),
  4726 => std_logic_vector'(x"000010ba"),
  4727 => std_logic_vector'(x"4e015401"),
  4728 => std_logic_vector'(x"4e2b5403"),
  4729 => std_logic_vector'(x"4e265403"),
  4730 => std_logic_vector'(x"4e7c5403"),
  4731 => std_logic_vector'(x"4e5e5403"),
  4732 => std_logic_vector'(x"04547e02"),
  4733 => std_logic_vector'(x"543d3d4e"),
  4734 => std_logic_vector'(x"543c4e03"),
  4735 => std_logic_vector'(x"3e3e4e04"),
  4736 => std_logic_vector'(x"3c4e0454"),
  4737 => std_logic_vector'(x"7202543c"),
  4738 => std_logic_vector'(x"545b0354"),
  4739 => std_logic_vector'(x"6f69055d"),
  4740 => std_logic_vector'(x"065d545b"),
  4741 => std_logic_vector'(x"74617473"),
  4742 => std_logic_vector'(x"4e047375"),
  4743 => std_logic_vector'(x"00543c75"),
  4744 => std_logic_vector'(x"6f0349d2"),
  4745 => std_logic_vector'(x"10be3370"),
  4746 => std_logic_vector'(x"2d540400"),
  4747 => std_logic_vector'(x"54044e3e"),
  4748 => std_logic_vector'(x"06523e2d"),
  4749 => std_logic_vector'(x"5b3e2d4e"),
  4750 => std_logic_vector'(x"4e085d54"),
  4751 => std_logic_vector'(x"6f693e2d"),
  4752 => std_logic_vector'(x"065d545b"),
  4753 => std_logic_vector'(x"524f495f"),
  4754 => std_logic_vector'(x"4a205f44"),
  4755 => std_logic_vector'(x"72706f03"),
  4756 => std_logic_vector'(x"000010c2"),
  4757 => std_logic_vector'(x"2b720300"),
  4758 => std_logic_vector'(x"72030031"),
  4759 => std_logic_vector'(x"4a4a312d"),
  4760 => std_logic_vector'(x"64706f03"),
  4761 => std_logic_vector'(x"000010c6"),
  4762 => std_logic_vector'(x"2b640300"),
  4763 => std_logic_vector'(x"64030031"),
  4764 => std_logic_vector'(x"4a5e312d"),
  4765 => std_logic_vector'(x"696b7306"),
  4766 => std_logic_vector'(x"00222e70"),
  4767 => std_logic_vector'(x"4a7210ca"),
  4768 => std_logic_vector'(x"6c612e04"),
  4769 => std_logic_vector'(x"10e80075"),
  4770 => std_logic_vector'(x"554c4104"),
  4771 => std_logic_vector'(x"003b0120"),
  4772 => std_logic_vector'(x"4a044a7e"),
  4773 => std_logic_vector'(x"00706f31"),
  4774 => std_logic_vector'(x"00001144"),
  4775 => std_logic_vector'(x"0000113a"),
  4776 => std_logic_vector'(x"00001130"),
  4777 => std_logic_vector'(x"0000107c"),
  4778 => std_logic_vector'(x"0000112a"),
  4779 => std_logic_vector'(x"73034a90"),
  4780 => std_logic_vector'(x"11486565"),
  4781 => std_logic_vector'(x"650c4aac"),
  4782 => std_logic_vector'(x"7269766e"),
  4783 => std_logic_vector'(x"656d6e6f"),
  4784 => std_logic_vector'(x"003f746e"),
  4785 => std_logic_vector'(x"4ab411b0"),
  4786 => std_logic_vector'(x"6c616608"),
  4787 => std_logic_vector'(x"656e6769"),
  4788 => std_logic_vector'(x"11b60064"),
  4789 => std_logic_vector'(x"66064ac6"),
  4790 => std_logic_vector'(x"74616f6c"),
  4791 => std_logic_vector'(x"11ba0073"),
  4792 => std_logic_vector'(x"73054ad4"),
  4793 => std_logic_vector'(x"3f656d61"),
  4794 => std_logic_vector'(x"4ae011be"),
  4795 => std_logic_vector'(x"6d6f6307"),
  4796 => std_logic_vector'(x"65726170"),
  4797 => std_logic_vector'(x"4aea11f6"),
  4798 => std_logic_vector'(x"616c6205"),
  4799 => std_logic_vector'(x"121c6b6e"),
  4800 => std_logic_vector'(x"2d094af6"),
  4801 => std_logic_vector'(x"69617274"),
  4802 => std_logic_vector'(x"676e696c"),
  4803 => std_logic_vector'(x"4b001222"),
  4804 => std_logic_vector'(x"61657306"),
  4805 => std_logic_vector'(x"00686372"),
  4806 => std_logic_vector'(x"4b0e123a"),
  4807 => std_logic_vector'(x"12843f01"),
  4808 => std_logic_vector'(x"28044b1a"),
  4809 => std_logic_vector'(x"0029732e"),
  4810 => std_logic_vector'(x"4b20128a"),
  4811 => std_logic_vector'(x"00732e02"),
  4812 => std_logic_vector'(x"4b2a129a"),
  4813 => std_logic_vector'(x"78656805"),
  4814 => std_logic_vector'(x"12ae2e32"),
  4815 => std_logic_vector'(x"64044b32"),
  4816 => std_logic_vector'(x"00706d75"),
  4817 => std_logic_vector'(x"4b3d12ca"),
  4818 => std_logic_vector'(x"4c455b06"),
  4819 => std_logic_vector'(x"005d4553"),
  4820 => std_logic_vector'(x"5b041350"),
  4821 => std_logic_vector'(x"065d4649"),
  4822 => std_logic_vector'(x"534c455b"),
  4823 => std_logic_vector'(x"5b065d45"),
  4824 => std_logic_vector'(x"4e454854"),
  4825 => std_logic_vector'(x"4b47005d"),
  4826 => std_logic_vector'(x"46495b04"),
  4827 => std_logic_vector'(x"13a4005d"),
  4828 => std_logic_vector'(x"5b064b67"),
  4829 => std_logic_vector'(x"4e454854"),
  4830 => std_logic_vector'(x"13ac005d"),
  4831 => std_logic_vector'(x"63074b70"),
  4832 => std_logic_vector'(x"69702d73"),
  4833 => std_logic_vector'(x"13ae6b63"),
  4834 => std_logic_vector'(x"63074b7c"),
  4835 => std_logic_vector'(x"6f722d73"),
  4836 => std_logic_vector'(x"13b26c6c"),
  4837 => std_logic_vector'(x"5b094b89"),
  4838 => std_logic_vector'(x"69666564"),
  4839 => std_logic_vector'(x"5d64656e"),
  4840 => std_logic_vector'(x"4b9513b6"),
  4841 => std_logic_vector'(x"6e755b0b"),
  4842 => std_logic_vector'(x"69666564"),
  4843 => std_logic_vector'(x"5d64656e"),
  4844 => std_logic_vector'(x"4ba213c4"),
  4845 => std_logic_vector'(x"6c617605"),
  4846 => std_logic_vector'(x"13ca6575"),
  4847 => std_logic_vector'(x"32064bb2"),
  4848 => std_logic_vector'(x"756c6176"),
  4849 => std_logic_vector'(x"13da0065"),
  4850 => std_logic_vector'(x"74024bbd"),
  4851 => std_logic_vector'(x"13ec006f"),
  4852 => std_logic_vector'(x"61084bc8"),
  4853 => std_logic_vector'(x"74726f62"),
  4854 => std_logic_vector'(x"0067736d"),
  4855 => std_logic_vector'(x"0000140a"),
  4856 => std_logic_vector'(x"00000000"),
  4857 => std_logic_vector'(x"28084bd0"),
  4858 => std_logic_vector'(x"726f6261"),
  4859 => std_logic_vector'(x"00292274"),
  4860 => std_logic_vector'(x"4be5140e"),
  4861 => std_logic_vector'(x"6f626106"),
  4862 => std_logic_vector'(x"00227472"),
  4863 => std_logic_vector'(x"4bf21422"),
  4864 => std_logic_vector'(x"69736303"),
  4865 => std_logic_vector'(x"4bfe142a"),
  4866 => std_logic_vector'(x"2d746105"),
  4867 => std_logic_vector'(x"14347978"),
  4868 => std_logic_vector'(x"70044c06"),
  4869 => std_logic_vector'(x"00656761"),
  4870 => std_logic_vector'(x"4c10144c"),
  4871 => std_logic_vector'(x"434f4c0a"),
  4872 => std_logic_vector'(x"4f574c41"),
  4873 => std_logic_vector'(x"00534452"),
  4874 => std_logic_vector'(x"4c1a145a"),
  4875 => std_logic_vector'(x"4255500b"),
  4876 => std_logic_vector'(x"5743494c"),
  4877 => std_logic_vector'(x"5344524f"),
  4878 => std_logic_vector'(x"4c2a145c"),
  4879 => std_logic_vector'(x"4e4f4409"),
  4880 => std_logic_vector'(x"524f5745"),
  4881 => std_logic_vector'(x"145e5344"),
  4882 => std_logic_vector'(x"63034c3a"),
  4883 => std_logic_vector'(x"1460212b"),
  4884 => std_logic_vector'(x"61074c48"),
  4885 => std_logic_vector'(x"68636464"),
  4886 => std_logic_vector'(x"146c7261"),
  4887 => std_logic_vector'(x"61064c50"),
  4888 => std_logic_vector'(x"6e657070"),
  4889 => std_logic_vector'(x"147c0064"),
  4890 => std_logic_vector'(x"65094c5c"),
  4891 => std_logic_vector'(x"61727478"),
  4892 => std_logic_vector'(x"48327463"),
  4893 => std_logic_vector'(x"4c681490"),
  4894 => std_logic_vector'(x"6373450b"),
  4895 => std_logic_vector'(x"54657061"),
  4896 => std_logic_vector'(x"656c6261"),
  4897 => std_logic_vector'(x"000014b8"),
  4898 => std_logic_vector'(x"64630807"),
  4899 => std_logic_vector'(x"68670c1b"),
  4900 => std_logic_vector'(x"0a6b6a69"),
  4901 => std_logic_vector'(x"706f0a6d"),
  4902 => std_logic_vector'(x"09730d22"),
  4903 => std_logic_vector'(x"78770b75"),
  4904 => std_logic_vector'(x"4c760079"),
  4905 => std_logic_vector'(x"4c524305"),
  4906 => std_logic_vector'(x"14bc2446"),
  4907 => std_logic_vector'(x"000a0d02"),
  4908 => std_logic_vector'(x"61094ca2"),
  4909 => std_logic_vector'(x"73456464"),
  4910 => std_logic_vector'(x"65706163"),
  4911 => std_logic_vector'(x"4cb014c0"),
  4912 => std_logic_vector'(x"72617007"),
  4913 => std_logic_vector'(x"225c6573"),
  4914 => std_logic_vector'(x"4cbe1546"),
  4915 => std_logic_vector'(x"6165720b"),
  4916 => std_logic_vector'(x"63734564"),
  4917 => std_logic_vector'(x"64657061"),
  4918 => std_logic_vector'(x"4ccb158e"),
  4919 => std_logic_vector'(x"225c5303"),
  4920 => std_logic_vector'(x"4cda15a8"),
  4921 => std_logic_vector'(x"66656405"),
  4922 => std_logic_vector'(x"15b67265"),
  4923 => std_logic_vector'(x"64064ce2"),
  4924 => std_logic_vector'(x"72656665"),
  4925 => std_logic_vector'(x"15c40040"),
  4926 => std_logic_vector'(x"64064cec"),
  4927 => std_logic_vector'(x"72656665"),
  4928 => std_logic_vector'(x"15ca0021"),
  4929 => std_logic_vector'(x"69024cf9"),
  4930 => std_logic_vector'(x"15d00073"),
  4931 => std_logic_vector'(x"61094d05"),
  4932 => std_logic_vector'(x"6f697463"),
  4933 => std_logic_vector'(x"666f2d6e"),
  4934 => std_logic_vector'(x"4d0c15e4"),
  4935 => std_logic_vector'(x"4c4f4805"),
  4936 => std_logic_vector'(x"15f85344"),
  4937 => std_logic_vector'(x"42074d1a"),
  4938 => std_logic_vector'(x"45464655"),
  4939 => std_logic_vector'(x"160c3a52"),
  4940 => std_logic_vector'(x"620f4d24"),
  4941 => std_logic_vector'(x"6e696765"),
  4942 => std_logic_vector'(x"7274732d"),
  4943 => std_logic_vector'(x"75746375"),
  4944 => std_logic_vector'(x"16126572"),
  4945 => std_logic_vector'(x"650d4d30"),
  4946 => std_logic_vector'(x"732d646e"),
  4947 => std_logic_vector'(x"63757274"),
  4948 => std_logic_vector'(x"65727574"),
  4949 => std_logic_vector'(x"4d441622"),
  4950 => std_logic_vector'(x"49462b06"),
  4951 => std_logic_vector'(x"00444c45"),
  4952 => std_logic_vector'(x"4d561628"),
  4953 => std_logic_vector'(x"69666307"),
  4954 => std_logic_vector'(x"3a646c65"),
  4955 => std_logic_vector'(x"4d621638"),
  4956 => std_logic_vector'(x"65696606"),
  4957 => std_logic_vector'(x"003a646c"),
  4958 => std_logic_vector'(x"4d6e1640"),
  4959 => std_logic_vector'(x"69666607"),
  4960 => std_logic_vector'(x"3a646c65"),
  4961 => std_logic_vector'(x"4d7a164a"),
  4962 => std_logic_vector'(x"6f6f6e04"),
  4963 => std_logic_vector'(x"16540070"),
  4964 => std_logic_vector'(x"6f034d86"),
  4965 => std_logic_vector'(x"16566666"),
  4966 => std_logic_vector'(x"6f024d90"),
  4967 => std_logic_vector'(x"165e006e"),
  4968 => std_logic_vector'(x"73044d98"),
  4969 => std_logic_vector'(x"00646565"),
  4970 => std_logic_vector'(x"00001666"),
  4971 => std_logic_vector'(x"7a92764b"),
  4972 => std_logic_vector'(x"73074da0"),
  4973 => std_logic_vector'(x"65737465"),
  4974 => std_logic_vector'(x"166a6465"),
  4975 => std_logic_vector'(x"72064db0"),
  4976 => std_logic_vector'(x"6f646e61"),
  4977 => std_logic_vector'(x"1676006d"),
  4978 => std_logic_vector'(x"72094dbc"),
  4979 => std_logic_vector'(x"72646e61"),
  4980 => std_logic_vector'(x"65676e61"),
  4981 => std_logic_vector'(x"4dc8169a"),
  4982 => std_logic_vector'(x"746f6e03"),
  4983 => std_logic_vector'(x"4dd616a2"),
  4984 => std_logic_vector'(x"74656d06"),
  4985 => std_logic_vector'(x"00646f68"),
  4986 => std_logic_vector'(x"4dde16a6"),
  4987 => std_logic_vector'(x"72617603"),
  4988 => std_logic_vector'(x"4dea16c2"),
  4989 => std_logic_vector'(x"616c6305"),
  4990 => std_logic_vector'(x"16d27373"),
  4991 => std_logic_vector'(x"65094df2"),
  4992 => std_logic_vector'(x"632d646e"),
  4993 => std_logic_vector'(x"7373616c"),
  4994 => std_logic_vector'(x"4dfc16d8"),
  4995 => std_logic_vector'(x"74763e03"),
  4996 => std_logic_vector'(x"4e0a1716"),
  4997 => std_logic_vector'(x"6e696204"),
  4998 => std_logic_vector'(x"17200064"),
  4999 => std_logic_vector'(x"64074e12"),
  5000 => std_logic_vector'(x"6e696665"),
  5001 => std_logic_vector'(x"17267365"),
  5002 => std_logic_vector'(x"61044e1c"),
  5003 => std_logic_vector'(x"0077656e"),
  5004 => std_logic_vector'(x"4e28172c"),
  5005 => std_logic_vector'(x"003a3a02"),
  5006 => std_logic_vector'(x"4e32173c"),
  5007 => std_logic_vector'(x"6a626f06"),
  5008 => std_logic_vector'(x"00746365"),
  5009 => std_logic_vector'(x"00001742"),
  5010 => std_logic_vector'(x"00000004"),
  5011 => std_logic_vector'(x"00000008"),
  5012 => std_logic_vector'(x"49054e3a"),
  5013 => std_logic_vector'(x"5455504e"),
  5014 => std_logic_vector'(x"4e501746"),
  5015 => std_logic_vector'(x"54554f06"),
  5016 => std_logic_vector'(x"00545550"),
  5017 => std_logic_vector'(x"4e5a174a"),
  5018 => std_logic_vector'(x"6e697007"),
  5019 => std_logic_vector'(x"65646f4d"),
  5020 => std_logic_vector'(x"4e66174e"),
  5021 => std_logic_vector'(x"6769640b"),
  5022 => std_logic_vector'(x"6c617469"),
  5023 => std_logic_vector'(x"64616552"),
  5024 => std_logic_vector'(x"4e721756"),
  5025 => std_logic_vector'(x"6769640c"),
  5026 => std_logic_vector'(x"6c617469"),
  5027 => std_logic_vector'(x"74697257"),
  5028 => std_logic_vector'(x"175a0065"),
  5029 => std_logic_vector'(x"74054e82"),
  5030 => std_logic_vector'(x"626f7268"),
  5031 => std_logic_vector'(x"4e94175e"),
  5032 => std_logic_vector'(x"006f6c02"),
  5033 => std_logic_vector'(x"4e9e1774"),
  5034 => std_logic_vector'(x"00696802"),
  5035 => std_logic_vector'(x"4ea6177c"),
  5036 => std_logic_vector'(x"534f4d04"),
  5037 => std_logic_vector'(x"17840049"),
  5038 => std_logic_vector'(x"4d044eae"),
  5039 => std_logic_vector'(x"004f5349"),
  5040 => std_logic_vector'(x"4eb81788"),
  5041 => std_logic_vector'(x"4b435303"),
  5042 => std_logic_vector'(x"4ec2178c"),
  5043 => std_logic_vector'(x"69627804"),
  5044 => std_logic_vector'(x"17900074"),
  5045 => std_logic_vector'(x"73044eca"),
  5046 => std_logic_vector'(x"00786970"),
  5047 => std_logic_vector'(x"4ed417a4"),
  5048 => std_logic_vector'(x"69707304"),
  5049 => std_logic_vector'(x"17dc003e"),
  5050 => std_logic_vector'(x"73084ede"),
  5051 => std_logic_vector'(x"692d6970"),
  5052 => std_logic_vector'(x"0074696e"),
  5053 => std_logic_vector'(x"4ee817e2"),
  5054 => std_logic_vector'(x"70733e04"),
  5055 => std_logic_vector'(x"17f00069"),
  5056 => std_logic_vector'(x"62074ef6"),
  5057 => std_logic_vector'(x"733e6b6c"),
  5058 => std_logic_vector'(x"18206970"),
  5059 => std_logic_vector'(x"66044f00"),
  5060 => std_logic_vector'(x"00716572"),
  5061 => std_logic_vector'(x"4f0c1838"),
  5062 => std_logic_vector'(x"6b6c6304"),
  5063 => std_logic_vector'(x"183e0040"),
  5064 => std_logic_vector'(x"74024f16"),
  5065 => std_logic_vector'(x"184e0075"),
  5066 => std_logic_vector'(x"6d034f20"),
  5067 => std_logic_vector'(x"18584073"),
  5068 => std_logic_vector'(x"75034f28"),
  5069 => std_logic_vector'(x"185e4073"),
  5070 => std_logic_vector'(x"6e034f30"),
  5071 => std_logic_vector'(x"186c4073"),
  5072 => std_logic_vector'(x"6d024f38"),
  5073 => std_logic_vector'(x"187a0073"),
  5074 => std_logic_vector'(x"6e034f40"),
  5075 => std_logic_vector'(x"18927765"),
  5076 => std_logic_vector'(x"6d207c0a"),
  5077 => std_logic_vector'(x"656b7261"),
  5078 => std_logic_vector'(x"007c2072"),
  5079 => std_logic_vector'(x"7c014f48"),
  5080 => std_logic_vector'(x"0000189a"),
  5081 => std_logic_vector'(x"0000189a"),
  5082 => std_logic_vector'(x"00004f5b"),
  5083 => std_logic_vector'(x"00004f48"),
  5084 => std_logic_vector'(x"55054f5c"),
  5085 => std_logic_vector'(x"73657244"),
  5086 => std_logic_vector'(x"0000189e"),
  5087 => std_logic_vector'(x"00071afd"),
  5088 => std_logic_vector'(x"4b56c380"),
  5089 => std_logic_vector'(x"00132f4a"),
  5090 => std_logic_vector'(x"e6c93315"),
  5091 => std_logic_vector'(x"63084f70"),
  5092 => std_logic_vector'(x"5f6c6c65"),
  5093 => std_logic_vector'(x"0062736d"),
  5094 => std_logic_vector'(x"4f8c18a2"),
  5095 => std_logic_vector'(x"3c647503"),
  5096 => std_logic_vector'(x"4f9a18b8"),
  5097 => std_logic_vector'(x"3c6e7503"),
  5098 => std_logic_vector'(x"4fa218d6"),
  5099 => std_logic_vector'(x"2d6e7503"),
  5100 => std_logic_vector'(x"4faa1928"),
  5101 => std_logic_vector'(x"2f326e03"),
  5102 => std_logic_vector'(x"4fb21990"),
  5103 => std_logic_vector'(x"2a647503"),
  5104 => std_logic_vector'(x"4fba19d2"),
  5105 => std_logic_vector'(x"73445505"),
  5106 => std_logic_vector'(x"1a5c6275"),
  5107 => std_logic_vector'(x"00038d7e"),
  5108 => std_logic_vector'(x"a69f85c0"),
  5109 => std_logic_vector'(x"00132f4a"),
  5110 => std_logic_vector'(x"e6c673f5"),
  5111 => std_logic_vector'(x"2e064fc2"),
  5112 => std_logic_vector'(x"75734455"),
  5113 => std_logic_vector'(x"1a600062"),
  5114 => std_logic_vector'(x"73445507"),
  5115 => std_logic_vector'(x"203a6275"),
  5116 => std_logic_vector'(x"2e064fdc"),
  5117 => std_logic_vector'(x"65724455"),
  5118 => std_logic_vector'(x"1a860073"),
  5119 => std_logic_vector'(x"72445507"),
  5120 => std_logic_vector'(x"203a7365"),
  5121 => std_logic_vector'(x"75034ff0"),
  5122 => std_logic_vector'(x"1aac2f64"),
  5123 => std_logic_vector'(x"65764f08"),
  5124 => std_logic_vector'(x"6f6c6672"),
  5125 => std_logic_vector'(x"50040077"),
  5126 => std_logic_vector'(x"40647503"),
  5127 => std_logic_vector'(x"50161b0e"),
  5128 => std_logic_vector'(x"43324908"),
  5129 => std_logic_vector'(x"4745525f"),
  5130 => std_logic_vector'(x"1b220053"),
  5131 => std_logic_vector'(x"6508501e"),
  5132 => std_logic_vector'(x"685f7272"),
  5133 => std_logic_vector'(x"00746c61"),
  5134 => std_logic_vector'(x"502c1b26"),
  5135 => std_logic_vector'(x"63326908"),
  5136 => std_logic_vector'(x"696e695f"),
  5137 => std_logic_vector'(x"1b2e0074"),
  5138 => std_logic_vector'(x"6907503a"),
  5139 => std_logic_vector'(x"735f6332"),
  5140 => std_logic_vector'(x"1b4a766c"),
  5141 => std_logic_vector'(x"69075048"),
  5142 => std_logic_vector'(x"775f6332"),
  5143 => std_logic_vector'(x"1b803172"),
  5144 => std_logic_vector'(x"69075054"),
  5145 => std_logic_vector'(x"725f6332"),
  5146 => std_logic_vector'(x"1bba3164"),
  5147 => std_logic_vector'(x"69065060"),
  5148 => std_logic_vector'(x"775f6332"),
  5149 => std_logic_vector'(x"1bf20072"),
  5150 => std_logic_vector'(x"6906506c"),
  5151 => std_logic_vector'(x"725f6332"),
  5152 => std_logic_vector'(x"1c4c0064"),
  5153 => std_logic_vector'(x"46085078"),
  5154 => std_logic_vector'(x"5f305152"),
  5155 => std_logic_vector'(x"00544e43"),
  5156 => std_logic_vector'(x"50841cc4"),
  5157 => std_logic_vector'(x"51524608"),
  5158 => std_logic_vector'(x"4e435f31"),
  5159 => std_logic_vector'(x"1cc80054"),
  5160 => std_logic_vector'(x"46085092"),
  5161 => std_logic_vector'(x"5f325152"),
  5162 => std_logic_vector'(x"00544e43"),
  5163 => std_logic_vector'(x"50a01ccc"),
  5164 => std_logic_vector'(x"54554f08"),
  5165 => std_logic_vector'(x"45525f30"),
  5166 => std_logic_vector'(x"1cd00047"),
  5167 => std_logic_vector'(x"4f0850ae"),
  5168 => std_logic_vector'(x"5f315455"),
  5169 => std_logic_vector'(x"00474552"),
  5170 => std_logic_vector'(x"50bc1cd4"),
  5171 => std_logic_vector'(x"54554f08"),
  5172 => std_logic_vector'(x"45525f32"),
  5173 => std_logic_vector'(x"1cd80047"),
  5174 => std_logic_vector'(x"4f0850ca"),
  5175 => std_logic_vector'(x"5f335455"),
  5176 => std_logic_vector'(x"00474552"),
  5177 => std_logic_vector'(x"50d81cdc"),
  5178 => std_logic_vector'(x"504e4908"),
  5179 => std_logic_vector'(x"45525f30"),
  5180 => std_logic_vector'(x"1ce00047"),
  5181 => std_logic_vector'(x"490850e6"),
  5182 => std_logic_vector'(x"5f31504e"),
  5183 => std_logic_vector'(x"00474552"),
  5184 => std_logic_vector'(x"50f41ce4"),
  5185 => std_logic_vector'(x"504e4908"),
  5186 => std_logic_vector'(x"45525f32"),
  5187 => std_logic_vector'(x"1ce80047"),
  5188 => std_logic_vector'(x"49085102"),
  5189 => std_logic_vector'(x"5f33504e"),
  5190 => std_logic_vector'(x"00474552"),
  5191 => std_logic_vector'(x"51101cec"),
  5192 => std_logic_vector'(x"4332490b"),
  5193 => std_logic_vector'(x"5355425f"),
  5194 => std_logic_vector'(x"4c45535f"),
  5195 => std_logic_vector'(x"511e1cf0"),
  5196 => std_logic_vector'(x"73756207"),
  5197 => std_logic_vector'(x"6c65735f"),
  5198 => std_logic_vector'(x"512e1cf4"),
  5199 => std_logic_vector'(x"43324907"),
  5200 => std_logic_vector'(x"58554d5f"),
  5201 => std_logic_vector'(x"513a1cfa"),
  5202 => std_logic_vector'(x"4332490d"),
  5203 => std_logic_vector'(x"58554d5f"),
  5204 => std_logic_vector'(x"3569535f"),
  5205 => std_logic_vector'(x"1cfe7837"),
  5206 => std_logic_vector'(x"490f5146"),
  5207 => std_logic_vector'(x"4d5f4332"),
  5208 => std_logic_vector'(x"415f5855"),
  5209 => std_logic_vector'(x"36344e44"),
  5210 => std_logic_vector'(x"1d023430"),
  5211 => std_logic_vector'(x"49085158"),
  5212 => std_logic_vector'(x"325f4332"),
  5213 => std_logic_vector'(x"00667562"),
  5214 => std_logic_vector'(x"00001d06"),
  5215 => std_logic_vector'(x"00000002"),
  5216 => std_logic_vector'(x"490a516c"),
  5217 => std_logic_vector'(x"695f4332"),
  5218 => std_logic_vector'(x"725f646e"),
  5219 => std_logic_vector'(x"1d0a0064"),
  5220 => std_logic_vector'(x"490a5180"),
  5221 => std_logic_vector'(x"695f4332"),
  5222 => std_logic_vector'(x"775f646e"),
  5223 => std_logic_vector'(x"1d140072"),
  5224 => std_logic_vector'(x"41075190"),
  5225 => std_logic_vector'(x"36344e44"),
  5226 => std_logic_vector'(x"1d2c3430"),
  5227 => std_logic_vector'(x"410a51a0"),
  5228 => std_logic_vector'(x"36344e44"),
  5229 => std_logic_vector'(x"725f3430"),
  5230 => std_logic_vector'(x"1d300064"),
  5231 => std_logic_vector'(x"410a51ac"),
  5232 => std_logic_vector'(x"36344e44"),
  5233 => std_logic_vector'(x"775f3430"),
  5234 => std_logic_vector'(x"1d360072"),
  5235 => std_logic_vector'(x"530551bc"),
  5236 => std_logic_vector'(x"78373569"),
  5237 => std_logic_vector'(x"51cc1d3c"),
  5238 => std_logic_vector'(x"3569530d"),
  5239 => std_logic_vector'(x"6f5f7837"),
  5240 => std_logic_vector'(x"6d5f646c"),
  5241 => std_logic_vector'(x"1d407875"),
  5242 => std_logic_vector'(x"00000000"),
  5243 => std_logic_vector'(x"530851d6"),
  5244 => std_logic_vector'(x"78373569"),
  5245 => std_logic_vector'(x"0072775f"),
  5246 => std_logic_vector'(x"51ec1d44"),
  5247 => std_logic_vector'(x"35695308"),
  5248 => std_logic_vector'(x"725f7837"),
  5249 => std_logic_vector'(x"1d4a0064"),
  5250 => std_logic_vector'(x"530851fa"),
  5251 => std_logic_vector'(x"46525f35"),
  5252 => std_logic_vector'(x"00514552"),
  5253 => std_logic_vector'(x"00001d50"),
  5254 => std_logic_vector'(x"00000000"),
  5255 => std_logic_vector'(x"00000000"),
  5256 => std_logic_vector'(x"53075208"),
  5257 => std_logic_vector'(x"44465f35"),
  5258 => std_logic_vector'(x"1d544f43"),
  5259 => std_logic_vector'(x"00000000"),
  5260 => std_logic_vector'(x"00000000"),
  5261 => std_logic_vector'(x"53055220"),
  5262 => std_logic_vector'(x"314e5f35"),
  5263 => std_logic_vector'(x"00001d58"),
  5264 => std_logic_vector'(x"00000000"),
  5265 => std_logic_vector'(x"53085234"),
  5266 => std_logic_vector'(x"53485f35"),
  5267 => std_logic_vector'(x"00564944"),
  5268 => std_logic_vector'(x"00001d5c"),
  5269 => std_logic_vector'(x"00000000"),
  5270 => std_logic_vector'(x"53085244"),
  5271 => std_logic_vector'(x"58465f35"),
  5272 => std_logic_vector'(x"004c4154"),
  5273 => std_logic_vector'(x"00001d60"),
  5274 => std_logic_vector'(x"00000000"),
  5275 => std_logic_vector'(x"310b5258"),
  5276 => std_logic_vector'(x"36453030"),
  5277 => std_logic_vector'(x"3c3c312a"),
  5278 => std_logic_vector'(x"1d643832"),
  5279 => std_logic_vector'(x"005f5e10"),
  5280 => std_logic_vector'(x"00000000"),
  5281 => std_logic_vector'(x"5308526c"),
  5282 => std_logic_vector'(x"44465f35"),
  5283 => std_logic_vector'(x"004c4f43"),
  5284 => std_logic_vector'(x"00001d68"),
  5285 => std_logic_vector'(x"00000001"),
  5286 => std_logic_vector'(x"21152080"),
  5287 => std_logic_vector'(x"53085284"),
  5288 => std_logic_vector'(x"44465f35"),
  5289 => std_logic_vector'(x"00484f43"),
  5290 => std_logic_vector'(x"00001d6c"),
  5291 => std_logic_vector'(x"00000001"),
  5292 => std_logic_vector'(x"51f55580"),
  5293 => std_logic_vector'(x"7308529c"),
  5294 => std_logic_vector'(x"73685f35"),
  5295 => std_logic_vector'(x"00737664"),
  5296 => std_logic_vector'(x"00001d70"),
  5297 => std_logic_vector'(x"0000000b"),
  5298 => std_logic_vector'(x"00000009"),
  5299 => std_logic_vector'(x"00000007"),
  5300 => std_logic_vector'(x"00000006"),
  5301 => std_logic_vector'(x"00000005"),
  5302 => std_logic_vector'(x"00000004"),
  5303 => std_logic_vector'(x"531052b4"),
  5304 => std_logic_vector'(x"78373569"),
  5305 => std_logic_vector'(x"6165725f"),
  5306 => std_logic_vector'(x"65735f64"),
  5307 => std_logic_vector'(x"00736774"),
  5308 => std_logic_vector'(x"52dc1d74"),
  5309 => std_logic_vector'(x"35695314"),
  5310 => std_logic_vector'(x"735f7837"),
  5311 => std_logic_vector'(x"725f6d69"),
  5312 => std_logic_vector'(x"5f646165"),
  5313 => std_logic_vector'(x"67746573"),
  5314 => std_logic_vector'(x"1dea0073"),
  5315 => std_logic_vector'(x"531052f2"),
  5316 => std_logic_vector'(x"78373569"),
  5317 => std_logic_vector'(x"6f68735f"),
  5318 => std_logic_vector'(x"65735f77"),
  5319 => std_logic_vector'(x"00736774"),
  5320 => std_logic_vector'(x"48071e0a"),
  5321 => std_logic_vector'(x"49445f53"),
  5322 => std_logic_vector'(x"4e033d56"),
  5323 => std_logic_vector'(x"46063d31"),
  5324 => std_logic_vector'(x"4c415458"),
  5325 => std_logic_vector'(x"4652063d"),
  5326 => std_logic_vector'(x"3d514552"),
  5327 => std_logic_vector'(x"43444605"),
  5328 => std_logic_vector'(x"46053d4f"),
  5329 => std_logic_vector'(x"3d54554f"),
  5330 => std_logic_vector'(x"5310530c"),
  5331 => std_logic_vector'(x"78373569"),
  5332 => std_logic_vector'(x"6c61635f"),
  5333 => std_logic_vector'(x"65735f63"),
  5334 => std_logic_vector'(x"00736774"),
  5335 => std_logic_vector'(x"53481e6e"),
  5336 => std_logic_vector'(x"35695311"),
  5337 => std_logic_vector'(x"775f7837"),
  5338 => std_logic_vector'(x"65746972"),
  5339 => std_logic_vector'(x"7465735f"),
  5340 => std_logic_vector'(x"1f407367"),
  5341 => std_logic_vector'(x"530c535e"),
  5342 => std_logic_vector'(x"78373569"),
  5343 => std_logic_vector'(x"7465535f"),
  5344 => std_logic_vector'(x"00717246"),
  5345 => std_logic_vector'(x"53741fca"),
  5346 => std_logic_vector'(x"534d460a"),
  5347 => std_logic_vector'(x"5f513431"),
  5348 => std_logic_vector'(x"00524441"),
  5349 => std_logic_vector'(x"53861fec"),
  5350 => std_logic_vector'(x"534d4609"),
  5351 => std_logic_vector'(x"5f513431"),
  5352 => std_logic_vector'(x"1ff07277"),
  5353 => std_logic_vector'(x"46095396"),
  5354 => std_logic_vector'(x"3431534d"),
  5355 => std_logic_vector'(x"64725f51"),
  5356 => std_logic_vector'(x"53a41ff6"),
  5357 => std_logic_vector'(x"34315307"),
  5358 => std_logic_vector'(x"3050435f"),
  5359 => std_logic_vector'(x"00001ffc"),
  5360 => std_logic_vector'(x"00000000"),
  5361 => std_logic_vector'(x"530653b2"),
  5362 => std_logic_vector'(x"4e5f3431"),
  5363 => std_logic_vector'(x"20000030"),
  5364 => std_logic_vector'(x"00000000"),
  5365 => std_logic_vector'(x"530653c4"),
  5366 => std_logic_vector'(x"4d5f3431"),
  5367 => std_logic_vector'(x"20040030"),
  5368 => std_logic_vector'(x"00000000"),
  5369 => std_logic_vector'(x"530753d4"),
  5370 => std_logic_vector'(x"505f3431"),
  5371 => std_logic_vector'(x"20087356"),
  5372 => std_logic_vector'(x"00000001"),
  5373 => std_logic_vector'(x"00000002"),
  5374 => std_logic_vector'(x"00000004"),
  5375 => std_logic_vector'(x"00000005"),
  5376 => std_logic_vector'(x"530653e4"),
  5377 => std_logic_vector'(x"505f3431"),
  5378 => std_logic_vector'(x"200c0030"),
  5379 => std_logic_vector'(x"00000000"),
  5380 => std_logic_vector'(x"53075400"),
  5381 => std_logic_vector'(x"505f3431"),
  5382 => std_logic_vector'(x"20105630"),
  5383 => std_logic_vector'(x"00000000"),
  5384 => std_logic_vector'(x"53085410"),
  5385 => std_logic_vector'(x"465f3431"),
  5386 => std_logic_vector'(x"004f4356"),
  5387 => std_logic_vector'(x"00002014"),
  5388 => std_logic_vector'(x"00000000"),
  5389 => std_logic_vector'(x"00000000"),
  5390 => std_logic_vector'(x"53085420"),
  5391 => std_logic_vector'(x"465f3431"),
  5392 => std_logic_vector'(x"00464552"),
  5393 => std_logic_vector'(x"00002018"),
  5394 => std_logic_vector'(x"00000000"),
  5395 => std_logic_vector'(x"00000000"),
  5396 => std_logic_vector'(x"53095438"),
  5397 => std_logic_vector'(x"465f3431"),
  5398 => std_logic_vector'(x"3054554f"),
  5399 => std_logic_vector'(x"5450201c"),
  5400 => std_logic_vector'(x"34315309"),
  5401 => std_logic_vector'(x"4356465f"),
  5402 => std_logic_vector'(x"20284c4f"),
  5403 => std_logic_vector'(x"00000000"),
  5404 => std_logic_vector'(x"743aa380"),
  5405 => std_logic_vector'(x"5309545e"),
  5406 => std_logic_vector'(x"465f3431"),
  5407 => std_logic_vector'(x"484f4356"),
  5408 => std_logic_vector'(x"0000202c"),
  5409 => std_logic_vector'(x"00000000"),
  5410 => std_logic_vector'(x"9af8da00"),
  5411 => std_logic_vector'(x"460f5474"),
  5412 => std_logic_vector'(x"3431534d"),
  5413 => std_logic_vector'(x"69735f51"),
  5414 => std_logic_vector'(x"65725f6d"),
  5415 => std_logic_vector'(x"20306461"),
  5416 => std_logic_vector'(x"3431530c"),
  5417 => std_logic_vector'(x"2a304d5f"),
  5418 => std_logic_vector'(x"38315e32"),
  5419 => std_logic_vector'(x"3153073d"),
  5420 => std_logic_vector'(x"304e5f34"),
  5421 => std_logic_vector'(x"31530a3d"),
  5422 => std_logic_vector'(x"52465f34"),
  5423 => std_logic_vector'(x"3d304645"),
  5424 => std_logic_vector'(x"4611548c"),
  5425 => std_logic_vector'(x"3431534d"),
  5426 => std_logic_vector'(x"65725f51"),
  5427 => std_logic_vector'(x"735f6461"),
  5428 => std_logic_vector'(x"73677465"),
  5429 => std_logic_vector'(x"530c207c"),
  5430 => std_logic_vector'(x"4d5f3431"),
  5431 => std_logic_vector'(x"5e322a30"),
  5432 => std_logic_vector'(x"073d3831"),
  5433 => std_logic_vector'(x"5f343153"),
  5434 => std_logic_vector'(x"0a3d304e"),
  5435 => std_logic_vector'(x"5f343153"),
  5436 => std_logic_vector'(x"46455246"),
  5437 => std_logic_vector'(x"54c03d30"),
  5438 => std_logic_vector'(x"534d4611"),
  5439 => std_logic_vector'(x"5f513431"),
  5440 => std_logic_vector'(x"636c6163"),
  5441 => std_logic_vector'(x"7465735f"),
  5442 => std_logic_vector'(x"21387367"),
  5443 => std_logic_vector'(x"756f4607"),
  5444 => std_logic_vector'(x"2021646e"),
  5445 => std_logic_vector'(x"63766605"),
  5446 => std_logic_vector'(x"66053d6f"),
  5447 => std_logic_vector'(x"3d666572"),
  5448 => std_logic_vector'(x"776f4c14"),
  5449 => std_logic_vector'(x"20207265"),
  5450 => std_logic_vector'(x"7369204d"),
  5451 => std_logic_vector'(x"6f6f7420"),
  5452 => std_logic_vector'(x"67696220"),
  5453 => std_logic_vector'(x"3d4d0220"),
  5454 => std_logic_vector'(x"461254f6"),
  5455 => std_logic_vector'(x"3431534d"),
  5456 => std_logic_vector'(x"72775f51"),
  5457 => std_logic_vector'(x"5f657469"),
  5458 => std_logic_vector'(x"67746573"),
  5459 => std_logic_vector'(x"22340073"),
  5460 => std_logic_vector'(x"460d5538"),
  5461 => std_logic_vector'(x"3431534d"),
  5462 => std_logic_vector'(x"65535f51"),
  5463 => std_logic_vector'(x"71724674"),
  5464 => std_logic_vector'(x"555022e0"),
  5465 => std_logic_vector'(x"6b6c430d"),
  5466 => std_logic_vector'(x"5f78744d"),
  5467 => std_logic_vector'(x"4f746553"),
  5468 => std_logic_vector'(x"22e87475"),
  5469 => std_logic_vector'(x"695f6e1f"),
  5470 => std_logic_vector'(x"756d206e"),
  5471 => std_logic_vector'(x"62207473"),
  5472 => std_logic_vector'(x"65622065"),
  5473 => std_logic_vector'(x"65657774"),
  5474 => std_logic_vector'(x"312d206e"),
  5475 => std_logic_vector'(x"646e6120"),
  5476 => std_logic_vector'(x"20353120"),
  5477 => std_logic_vector'(x"6f5f6e1f"),
  5478 => std_logic_vector'(x"6d207475"),
  5479 => std_logic_vector'(x"20747375"),
  5480 => std_logic_vector'(x"62206562"),
  5481 => std_logic_vector'(x"65777465"),
  5482 => std_logic_vector'(x"30206e65"),
  5483 => std_logic_vector'(x"646e6120"),
  5484 => std_logic_vector'(x"20353120"),
  5485 => std_logic_vector'(x"45075562"),
  5486 => std_logic_vector'(x"625f4955"),
  5487 => std_logic_vector'(x"23986675"),
  5488 => std_logic_vector'(x"00000000"),
  5489 => std_logic_vector'(x"00000000"),
  5490 => std_logic_vector'(x"55b40000"),
  5491 => std_logic_vector'(x"32544107"),
  5492 => std_logic_vector'(x"43414d34"),
  5493 => std_logic_vector'(x"55ca239c"),
  5494 => std_logic_vector'(x"3254410f"),
  5495 => std_logic_vector'(x"43414d34"),
  5496 => std_logic_vector'(x"6332695f"),
  5497 => std_logic_vector'(x"6c65735f"),
  5498 => std_logic_vector'(x"55d623a0"),
  5499 => std_logic_vector'(x"49554508"),
  5500 => std_logic_vector'(x"6165725f"),
  5501 => std_logic_vector'(x"23a40064"),
  5502 => std_logic_vector'(x"2e0855ea"),
  5503 => std_logic_vector'(x"65747962"),
  5504 => std_logic_vector'(x"00667562"),
  5505 => std_logic_vector'(x"55f823be"),
  5506 => std_logic_vector'(x"4346410d"),
  5507 => std_logic_vector'(x"32695f4b"),
  5508 => std_logic_vector'(x"6e695f63"),
  5509 => std_logic_vector'(x"23dc7469"),
  5510 => std_logic_vector'(x"00000000"),
  5511 => std_logic_vector'(x"00000000"),
  5512 => std_logic_vector'(x"00000000"),
  5513 => std_logic_vector'(x"00000000"),
  5514 => std_logic_vector'(x"00000000"),
  5515 => std_logic_vector'(x"00000000"),
  5516 => std_logic_vector'(x"00000000"),
  5517 => std_logic_vector'(x"00000000"),
  5518 => std_logic_vector'(x"00000000"),
  5519 => std_logic_vector'(x"00000000"),
  5520 => std_logic_vector'(x"00000000"),
  5521 => std_logic_vector'(x"00000000"),
  5522 => std_logic_vector'(x"00000000"),
  5523 => std_logic_vector'(x"00000000"),
  5524 => std_logic_vector'(x"00000000"),
  5525 => std_logic_vector'(x"00000000"),
  5526 => std_logic_vector'(x"00000000"),
  5527 => std_logic_vector'(x"00000000"),
  5528 => std_logic_vector'(x"00000000"),
  5529 => std_logic_vector'(x"00000000"),
  5530 => std_logic_vector'(x"00000000"),
  5531 => std_logic_vector'(x"00000000"),
  5532 => std_logic_vector'(x"00000000"),
  5533 => std_logic_vector'(x"00000000"),
  5534 => std_logic_vector'(x"00000000"),
  5535 => std_logic_vector'(x"00000000"),
  5536 => std_logic_vector'(x"00000000"),
  5537 => std_logic_vector'(x"00000000"),
  5538 => std_logic_vector'(x"00000000"),
  5539 => std_logic_vector'(x"00000000"),
  5540 => std_logic_vector'(x"00000000"),
  5541 => std_logic_vector'(x"00000000"),
  5542 => std_logic_vector'(x"00000000"),
  5543 => std_logic_vector'(x"00000000"),
  5544 => std_logic_vector'(x"00000000"),
  5545 => std_logic_vector'(x"00000000"),
  5546 => std_logic_vector'(x"00000000"),
  5547 => std_logic_vector'(x"00000000"),
  5548 => std_logic_vector'(x"00000000"),
  5549 => std_logic_vector'(x"00000000"),
  5550 => std_logic_vector'(x"00000000"),
  5551 => std_logic_vector'(x"00000000"),
  5552 => std_logic_vector'(x"00000000"),
  5553 => std_logic_vector'(x"00000000"),
  5554 => std_logic_vector'(x"00000000"),
  5555 => std_logic_vector'(x"00000000"),
  5556 => std_logic_vector'(x"00000000"),
  5557 => std_logic_vector'(x"00000000"),
  5558 => std_logic_vector'(x"00000000"),
  5559 => std_logic_vector'(x"00000000"),
  5560 => std_logic_vector'(x"00000000"),
  5561 => std_logic_vector'(x"00000000"),
  5562 => std_logic_vector'(x"00000000"),
  5563 => std_logic_vector'(x"00000000"),
  5564 => std_logic_vector'(x"00000000"),
  5565 => std_logic_vector'(x"00000000"),
  5566 => std_logic_vector'(x"00000000"),
  5567 => std_logic_vector'(x"00000000"),
  5568 => std_logic_vector'(x"00000000"),
  5569 => std_logic_vector'(x"00000000"),
  5570 => std_logic_vector'(x"00000000"),
  5571 => std_logic_vector'(x"00000000"),
  5572 => std_logic_vector'(x"00000000"),
  5573 => std_logic_vector'(x"00000000"),
  5574 => std_logic_vector'(x"00000000"),
  5575 => std_logic_vector'(x"00000000"),
  5576 => std_logic_vector'(x"00000000"),
  5577 => std_logic_vector'(x"00000000"),
  5578 => std_logic_vector'(x"00000000"),
  5579 => std_logic_vector'(x"00000000"),
  5580 => std_logic_vector'(x"00000000"),
  5581 => std_logic_vector'(x"00000000"),
  5582 => std_logic_vector'(x"00000000"),
  5583 => std_logic_vector'(x"00000000"),
  5584 => std_logic_vector'(x"00000000"),
  5585 => std_logic_vector'(x"00000000"),
  5586 => std_logic_vector'(x"00000000"),
  5587 => std_logic_vector'(x"00000000"),
  5588 => std_logic_vector'(x"00000000"),
  5589 => std_logic_vector'(x"00000000"),
  5590 => std_logic_vector'(x"00000000"),
  5591 => std_logic_vector'(x"00000000"),
  5592 => std_logic_vector'(x"00000000"),
  5593 => std_logic_vector'(x"00000000"),
  5594 => std_logic_vector'(x"00000000"),
  5595 => std_logic_vector'(x"00000000"),
  5596 => std_logic_vector'(x"00000000"),
  5597 => std_logic_vector'(x"00000000"),
  5598 => std_logic_vector'(x"00000000"),
  5599 => std_logic_vector'(x"00000000"),
  5600 => std_logic_vector'(x"00000000"),
  5601 => std_logic_vector'(x"00000000"),
  5602 => std_logic_vector'(x"00000000"),
  5603 => std_logic_vector'(x"00000000"),
  5604 => std_logic_vector'(x"00000000"),
  5605 => std_logic_vector'(x"00000000"),
  5606 => std_logic_vector'(x"00000000"),
  5607 => std_logic_vector'(x"00000000"),
  5608 => std_logic_vector'(x"00000000"),
  5609 => std_logic_vector'(x"00000000"),
  5610 => std_logic_vector'(x"00000000"),
  5611 => std_logic_vector'(x"00000000"),
  5612 => std_logic_vector'(x"00000000"),
  5613 => std_logic_vector'(x"00000000"),
  5614 => std_logic_vector'(x"00000000"),
  5615 => std_logic_vector'(x"00000000"),
  5616 => std_logic_vector'(x"00000000"),
  5617 => std_logic_vector'(x"00000000"),
  5618 => std_logic_vector'(x"00000000"),
  5619 => std_logic_vector'(x"00000000"),
  5620 => std_logic_vector'(x"00000000"),
  5621 => std_logic_vector'(x"00000000"),
  5622 => std_logic_vector'(x"00000000"),
  5623 => std_logic_vector'(x"00000000"),
  5624 => std_logic_vector'(x"00000000"),
  5625 => std_logic_vector'(x"00000000"),
  5626 => std_logic_vector'(x"00000000"),
  5627 => std_logic_vector'(x"00000000"),
  5628 => std_logic_vector'(x"00000000"),
  5629 => std_logic_vector'(x"00000000"),
  5630 => std_logic_vector'(x"00000000"),
  5631 => std_logic_vector'(x"00000000"),
  5632 => std_logic_vector'(x"00000000"),
  5633 => std_logic_vector'(x"00000000"),
  5634 => std_logic_vector'(x"00000000"),
  5635 => std_logic_vector'(x"00000000"),
  5636 => std_logic_vector'(x"00000000"),
  5637 => std_logic_vector'(x"00000000"),
  5638 => std_logic_vector'(x"00000000"),
  5639 => std_logic_vector'(x"00000000"),
  5640 => std_logic_vector'(x"00000000"),
  5641 => std_logic_vector'(x"00000000"),
  5642 => std_logic_vector'(x"00000000"),
  5643 => std_logic_vector'(x"00000000"),
  5644 => std_logic_vector'(x"00000000"),
  5645 => std_logic_vector'(x"00000000"),
  5646 => std_logic_vector'(x"00000000"),
  5647 => std_logic_vector'(x"00000000"),
  5648 => std_logic_vector'(x"00000000"),
  5649 => std_logic_vector'(x"00000000"),
  5650 => std_logic_vector'(x"00000000"),
  5651 => std_logic_vector'(x"00000000"),
  5652 => std_logic_vector'(x"00000000"),
  5653 => std_logic_vector'(x"00000000"),
  5654 => std_logic_vector'(x"00000000"),
  5655 => std_logic_vector'(x"00000000"),
  5656 => std_logic_vector'(x"00000000"),
  5657 => std_logic_vector'(x"00000000"),
  5658 => std_logic_vector'(x"00000000"),
  5659 => std_logic_vector'(x"00000000"),
  5660 => std_logic_vector'(x"00000000"),
  5661 => std_logic_vector'(x"00000000"),
  5662 => std_logic_vector'(x"00000000"),
  5663 => std_logic_vector'(x"00000000"),
  5664 => std_logic_vector'(x"00000000"),
  5665 => std_logic_vector'(x"00000000"),
  5666 => std_logic_vector'(x"00000000"),
  5667 => std_logic_vector'(x"00000000"),
  5668 => std_logic_vector'(x"00000000"),
  5669 => std_logic_vector'(x"00000000"),
  5670 => std_logic_vector'(x"00000000"),
  5671 => std_logic_vector'(x"00000000"),
  5672 => std_logic_vector'(x"00000000"),
  5673 => std_logic_vector'(x"00000000"),
  5674 => std_logic_vector'(x"00000000"),
  5675 => std_logic_vector'(x"00000000"),
  5676 => std_logic_vector'(x"00000000"),
  5677 => std_logic_vector'(x"00000000"),
  5678 => std_logic_vector'(x"00000000"),
  5679 => std_logic_vector'(x"00000000"),
  5680 => std_logic_vector'(x"00000000"),
  5681 => std_logic_vector'(x"00000000"),
  5682 => std_logic_vector'(x"00000000"),
  5683 => std_logic_vector'(x"00000000"),
  5684 => std_logic_vector'(x"00000000"),
  5685 => std_logic_vector'(x"00000000"),
  5686 => std_logic_vector'(x"00000000"),
  5687 => std_logic_vector'(x"00000000"),
  5688 => std_logic_vector'(x"00000000"),
  5689 => std_logic_vector'(x"00000000"),
  5690 => std_logic_vector'(x"00000000"),
  5691 => std_logic_vector'(x"00000000"),
  5692 => std_logic_vector'(x"00000000"),
  5693 => std_logic_vector'(x"00000000"),
  5694 => std_logic_vector'(x"00000000"),
  5695 => std_logic_vector'(x"00000000"),
  5696 => std_logic_vector'(x"00000000"),
  5697 => std_logic_vector'(x"00000000"),
  5698 => std_logic_vector'(x"00000000"),
  5699 => std_logic_vector'(x"00000000"),
  5700 => std_logic_vector'(x"00000000"),
  5701 => std_logic_vector'(x"00000000"),
  5702 => std_logic_vector'(x"00000000"),
  5703 => std_logic_vector'(x"00000000"),
  5704 => std_logic_vector'(x"00000000"),
  5705 => std_logic_vector'(x"00000000"),
  5706 => std_logic_vector'(x"00000000"),
  5707 => std_logic_vector'(x"00000000"),
  5708 => std_logic_vector'(x"00000000"),
  5709 => std_logic_vector'(x"00000000"),
  5710 => std_logic_vector'(x"00000000"),
  5711 => std_logic_vector'(x"00000000"),
  5712 => std_logic_vector'(x"00000000"),
  5713 => std_logic_vector'(x"00000000"),
  5714 => std_logic_vector'(x"00000000"),
  5715 => std_logic_vector'(x"00000000"),
  5716 => std_logic_vector'(x"00000000"),
  5717 => std_logic_vector'(x"00000000"),
  5718 => std_logic_vector'(x"00000000"),
  5719 => std_logic_vector'(x"00000000"),
  5720 => std_logic_vector'(x"00000000"),
  5721 => std_logic_vector'(x"00000000"),
  5722 => std_logic_vector'(x"00000000"),
  5723 => std_logic_vector'(x"00000000"),
  5724 => std_logic_vector'(x"00000000"),
  5725 => std_logic_vector'(x"00000000"),
  5726 => std_logic_vector'(x"00000000"),
  5727 => std_logic_vector'(x"00000000"),
  5728 => std_logic_vector'(x"00000000"),
  5729 => std_logic_vector'(x"00000000"),
  5730 => std_logic_vector'(x"00000000"),
  5731 => std_logic_vector'(x"00000000"),
  5732 => std_logic_vector'(x"00000000"),
  5733 => std_logic_vector'(x"00000000"),
  5734 => std_logic_vector'(x"00000000"),
  5735 => std_logic_vector'(x"00000000"),
  5736 => std_logic_vector'(x"00000000"),
  5737 => std_logic_vector'(x"00000000"),
  5738 => std_logic_vector'(x"00000000"),
  5739 => std_logic_vector'(x"00000000"),
  5740 => std_logic_vector'(x"00000000"),
  5741 => std_logic_vector'(x"00000000"),
  5742 => std_logic_vector'(x"00000000"),
  5743 => std_logic_vector'(x"00000000"),
  5744 => std_logic_vector'(x"00000000"),
  5745 => std_logic_vector'(x"00000000"),
  5746 => std_logic_vector'(x"00000000"),
  5747 => std_logic_vector'(x"00000000"),
  5748 => std_logic_vector'(x"00000000"),
  5749 => std_logic_vector'(x"00000000"),
  5750 => std_logic_vector'(x"00000000"),
  5751 => std_logic_vector'(x"00000000"),
  5752 => std_logic_vector'(x"00000000"),
  5753 => std_logic_vector'(x"00000000"),
  5754 => std_logic_vector'(x"00000000"),
  5755 => std_logic_vector'(x"00000000"),
  5756 => std_logic_vector'(x"00000000"),
  5757 => std_logic_vector'(x"00000000"),
  5758 => std_logic_vector'(x"00000000"),
  5759 => std_logic_vector'(x"00000000"),
  5760 => std_logic_vector'(x"00000000"),
  5761 => std_logic_vector'(x"00000000"),
  5762 => std_logic_vector'(x"00000000"),
  5763 => std_logic_vector'(x"00000000"),
  5764 => std_logic_vector'(x"00000000"),
  5765 => std_logic_vector'(x"00000000"),
  5766 => std_logic_vector'(x"00000000"),
  5767 => std_logic_vector'(x"00000000"),
  5768 => std_logic_vector'(x"00000000"),
  5769 => std_logic_vector'(x"00000000"),
  5770 => std_logic_vector'(x"00000000"),
  5771 => std_logic_vector'(x"00000000"),
  5772 => std_logic_vector'(x"00000000"),
  5773 => std_logic_vector'(x"00000000"),
  5774 => std_logic_vector'(x"00000000"),
  5775 => std_logic_vector'(x"00000000"),
  5776 => std_logic_vector'(x"00000000"),
  5777 => std_logic_vector'(x"00000000"),
  5778 => std_logic_vector'(x"00000000"),
  5779 => std_logic_vector'(x"00000000"),
  5780 => std_logic_vector'(x"00000000"),
  5781 => std_logic_vector'(x"00000000"),
  5782 => std_logic_vector'(x"00000000"),
  5783 => std_logic_vector'(x"00000000"),
  5784 => std_logic_vector'(x"00000000"),
  5785 => std_logic_vector'(x"00000000"),
  5786 => std_logic_vector'(x"00000000"),
  5787 => std_logic_vector'(x"00000000"),
  5788 => std_logic_vector'(x"00000000"),
  5789 => std_logic_vector'(x"00000000"),
  5790 => std_logic_vector'(x"00000000"),
  5791 => std_logic_vector'(x"00000000"),
  5792 => std_logic_vector'(x"00000000"),
  5793 => std_logic_vector'(x"00000000"),
  5794 => std_logic_vector'(x"00000000"),
  5795 => std_logic_vector'(x"00000000"),
  5796 => std_logic_vector'(x"00000000"),
  5797 => std_logic_vector'(x"00000000"),
  5798 => std_logic_vector'(x"00000000"),
  5799 => std_logic_vector'(x"00000000"),
  5800 => std_logic_vector'(x"00000000"),
  5801 => std_logic_vector'(x"00000000"),
  5802 => std_logic_vector'(x"00000000"),
  5803 => std_logic_vector'(x"00000000"),
  5804 => std_logic_vector'(x"00000000"),
  5805 => std_logic_vector'(x"00000000"),
  5806 => std_logic_vector'(x"00000000"),
  5807 => std_logic_vector'(x"00000000"),
  5808 => std_logic_vector'(x"00000000"),
  5809 => std_logic_vector'(x"00000000"),
  5810 => std_logic_vector'(x"00000000"),
  5811 => std_logic_vector'(x"00000000"),
  5812 => std_logic_vector'(x"00000000"),
  5813 => std_logic_vector'(x"00000000"),
  5814 => std_logic_vector'(x"00000000"),
  5815 => std_logic_vector'(x"00000000"),
  5816 => std_logic_vector'(x"00000000"),
  5817 => std_logic_vector'(x"00000000"),
  5818 => std_logic_vector'(x"00000000"),
  5819 => std_logic_vector'(x"00000000"),
  5820 => std_logic_vector'(x"00000000"),
  5821 => std_logic_vector'(x"00000000"),
  5822 => std_logic_vector'(x"00000000"),
  5823 => std_logic_vector'(x"00000000"),
  5824 => std_logic_vector'(x"00000000"),
  5825 => std_logic_vector'(x"00000000"),
  5826 => std_logic_vector'(x"00000000"),
  5827 => std_logic_vector'(x"00000000"),
  5828 => std_logic_vector'(x"00000000"),
  5829 => std_logic_vector'(x"00000000"),
  5830 => std_logic_vector'(x"00000000"),
  5831 => std_logic_vector'(x"00000000"),
  5832 => std_logic_vector'(x"00000000"),
  5833 => std_logic_vector'(x"00000000"),
  5834 => std_logic_vector'(x"00000000"),
  5835 => std_logic_vector'(x"00000000"),
  5836 => std_logic_vector'(x"00000000"),
  5837 => std_logic_vector'(x"00000000"),
  5838 => std_logic_vector'(x"00000000"),
  5839 => std_logic_vector'(x"00000000"),
  5840 => std_logic_vector'(x"00000000"),
  5841 => std_logic_vector'(x"00000000"),
  5842 => std_logic_vector'(x"00000000"),
  5843 => std_logic_vector'(x"00000000"),
  5844 => std_logic_vector'(x"00000000"),
  5845 => std_logic_vector'(x"00000000"),
  5846 => std_logic_vector'(x"00000000"),
  5847 => std_logic_vector'(x"00000000"),
  5848 => std_logic_vector'(x"00000000"),
  5849 => std_logic_vector'(x"00000000"),
  5850 => std_logic_vector'(x"00000000"),
  5851 => std_logic_vector'(x"00000000"),
  5852 => std_logic_vector'(x"00000000"),
  5853 => std_logic_vector'(x"00000000"),
  5854 => std_logic_vector'(x"00000000"),
  5855 => std_logic_vector'(x"00000000"),
  5856 => std_logic_vector'(x"00000000"),
  5857 => std_logic_vector'(x"00000000"),
  5858 => std_logic_vector'(x"00000000"),
  5859 => std_logic_vector'(x"00000000"),
  5860 => std_logic_vector'(x"00000000"),
  5861 => std_logic_vector'(x"00000000"),
  5862 => std_logic_vector'(x"00000000"),
  5863 => std_logic_vector'(x"00000000"),
  5864 => std_logic_vector'(x"00000000"),
  5865 => std_logic_vector'(x"00000000"),
  5866 => std_logic_vector'(x"00000000"),
  5867 => std_logic_vector'(x"00000000"),
  5868 => std_logic_vector'(x"00000000"),
  5869 => std_logic_vector'(x"00000000"),
  5870 => std_logic_vector'(x"00000000"),
  5871 => std_logic_vector'(x"00000000"),
  5872 => std_logic_vector'(x"00000000"),
  5873 => std_logic_vector'(x"00000000"),
  5874 => std_logic_vector'(x"00000000"),
  5875 => std_logic_vector'(x"00000000"),
  5876 => std_logic_vector'(x"00000000"),
  5877 => std_logic_vector'(x"00000000"),
  5878 => std_logic_vector'(x"00000000"),
  5879 => std_logic_vector'(x"00000000"),
  5880 => std_logic_vector'(x"00000000"),
  5881 => std_logic_vector'(x"00000000"),
  5882 => std_logic_vector'(x"00000000"),
  5883 => std_logic_vector'(x"00000000"),
  5884 => std_logic_vector'(x"00000000"),
  5885 => std_logic_vector'(x"00000000"),
  5886 => std_logic_vector'(x"00000000"),
  5887 => std_logic_vector'(x"00000000"),
  5888 => std_logic_vector'(x"00000000"),
  5889 => std_logic_vector'(x"00000000"),
  5890 => std_logic_vector'(x"00000000"),
  5891 => std_logic_vector'(x"00000000"),
  5892 => std_logic_vector'(x"00000000"),
  5893 => std_logic_vector'(x"00000000"),
  5894 => std_logic_vector'(x"00000000"),
  5895 => std_logic_vector'(x"00000000"),
  5896 => std_logic_vector'(x"00000000"),
  5897 => std_logic_vector'(x"00000000"),
  5898 => std_logic_vector'(x"00000000"),
  5899 => std_logic_vector'(x"00000000"),
  5900 => std_logic_vector'(x"00000000"),
  5901 => std_logic_vector'(x"00000000"),
  5902 => std_logic_vector'(x"00000000"),
  5903 => std_logic_vector'(x"00000000"),
  5904 => std_logic_vector'(x"00000000"),
  5905 => std_logic_vector'(x"00000000"),
  5906 => std_logic_vector'(x"00000000"),
  5907 => std_logic_vector'(x"00000000"),
  5908 => std_logic_vector'(x"00000000"),
  5909 => std_logic_vector'(x"00000000"),
  5910 => std_logic_vector'(x"00000000"),
  5911 => std_logic_vector'(x"00000000"),
  5912 => std_logic_vector'(x"00000000"),
  5913 => std_logic_vector'(x"00000000"),
  5914 => std_logic_vector'(x"00000000"),
  5915 => std_logic_vector'(x"00000000"),
  5916 => std_logic_vector'(x"00000000"),
  5917 => std_logic_vector'(x"00000000"),
  5918 => std_logic_vector'(x"00000000"),
  5919 => std_logic_vector'(x"00000000"),
  5920 => std_logic_vector'(x"00000000"),
  5921 => std_logic_vector'(x"00000000"),
  5922 => std_logic_vector'(x"00000000"),
  5923 => std_logic_vector'(x"00000000"),
  5924 => std_logic_vector'(x"00000000"),
  5925 => std_logic_vector'(x"00000000"),
  5926 => std_logic_vector'(x"00000000"),
  5927 => std_logic_vector'(x"00000000"),
  5928 => std_logic_vector'(x"00000000"),
  5929 => std_logic_vector'(x"00000000"),
  5930 => std_logic_vector'(x"00000000"),
  5931 => std_logic_vector'(x"00000000"),
  5932 => std_logic_vector'(x"00000000"),
  5933 => std_logic_vector'(x"00000000"),
  5934 => std_logic_vector'(x"00000000"),
  5935 => std_logic_vector'(x"00000000"),
  5936 => std_logic_vector'(x"00000000"),
  5937 => std_logic_vector'(x"00000000"),
  5938 => std_logic_vector'(x"00000000"),
  5939 => std_logic_vector'(x"00000000"),
  5940 => std_logic_vector'(x"00000000"),
  5941 => std_logic_vector'(x"00000000"),
  5942 => std_logic_vector'(x"00000000"),
  5943 => std_logic_vector'(x"00000000"),
  5944 => std_logic_vector'(x"00000000"),
  5945 => std_logic_vector'(x"00000000"),
  5946 => std_logic_vector'(x"00000000"),
  5947 => std_logic_vector'(x"00000000"),
  5948 => std_logic_vector'(x"00000000"),
  5949 => std_logic_vector'(x"00000000"),
  5950 => std_logic_vector'(x"00000000"),
  5951 => std_logic_vector'(x"00000000"),
  5952 => std_logic_vector'(x"00000000"),
  5953 => std_logic_vector'(x"00000000"),
  5954 => std_logic_vector'(x"00000000"),
  5955 => std_logic_vector'(x"00000000"),
  5956 => std_logic_vector'(x"00000000"),
  5957 => std_logic_vector'(x"00000000"),
  5958 => std_logic_vector'(x"00000000"),
  5959 => std_logic_vector'(x"00000000"),
  5960 => std_logic_vector'(x"00000000"),
  5961 => std_logic_vector'(x"00000000"),
  5962 => std_logic_vector'(x"00000000"),
  5963 => std_logic_vector'(x"00000000"),
  5964 => std_logic_vector'(x"00000000"),
  5965 => std_logic_vector'(x"00000000"),
  5966 => std_logic_vector'(x"00000000"),
  5967 => std_logic_vector'(x"00000000"),
  5968 => std_logic_vector'(x"00000000"),
  5969 => std_logic_vector'(x"00000000"),
  5970 => std_logic_vector'(x"00000000"),
  5971 => std_logic_vector'(x"00000000"),
  5972 => std_logic_vector'(x"00000000"),
  5973 => std_logic_vector'(x"00000000"),
  5974 => std_logic_vector'(x"00000000"),
  5975 => std_logic_vector'(x"00000000"),
  5976 => std_logic_vector'(x"00000000"),
  5977 => std_logic_vector'(x"00000000"),
  5978 => std_logic_vector'(x"00000000"),
  5979 => std_logic_vector'(x"00000000"),
  5980 => std_logic_vector'(x"00000000"),
  5981 => std_logic_vector'(x"00000000"),
  5982 => std_logic_vector'(x"00000000"),
  5983 => std_logic_vector'(x"00000000"),
  5984 => std_logic_vector'(x"00000000"),
  5985 => std_logic_vector'(x"00000000"),
  5986 => std_logic_vector'(x"00000000"),
  5987 => std_logic_vector'(x"00000000"),
  5988 => std_logic_vector'(x"00000000"),
  5989 => std_logic_vector'(x"00000000"),
  5990 => std_logic_vector'(x"00000000"),
  5991 => std_logic_vector'(x"00000000"),
  5992 => std_logic_vector'(x"00000000"),
  5993 => std_logic_vector'(x"00000000"),
  5994 => std_logic_vector'(x"00000000"),
  5995 => std_logic_vector'(x"00000000"),
  5996 => std_logic_vector'(x"00000000"),
  5997 => std_logic_vector'(x"00000000"),
  5998 => std_logic_vector'(x"00000000"),
  5999 => std_logic_vector'(x"00000000"),
  6000 => std_logic_vector'(x"00000000"),
  6001 => std_logic_vector'(x"00000000"),
  6002 => std_logic_vector'(x"00000000"),
  6003 => std_logic_vector'(x"00000000"),
  6004 => std_logic_vector'(x"00000000"),
  6005 => std_logic_vector'(x"00000000"),
  6006 => std_logic_vector'(x"00000000"),
  6007 => std_logic_vector'(x"00000000"),
  6008 => std_logic_vector'(x"00000000"),
  6009 => std_logic_vector'(x"00000000"),
  6010 => std_logic_vector'(x"00000000"),
  6011 => std_logic_vector'(x"00000000"),
  6012 => std_logic_vector'(x"00000000"),
  6013 => std_logic_vector'(x"00000000"),
  6014 => std_logic_vector'(x"00000000"),
  6015 => std_logic_vector'(x"00000000"),
  6016 => std_logic_vector'(x"00000000"),
  6017 => std_logic_vector'(x"00000000"),
  6018 => std_logic_vector'(x"00000000"),
  6019 => std_logic_vector'(x"00000000"),
  6020 => std_logic_vector'(x"00000000"),
  6021 => std_logic_vector'(x"00000000"),
  6022 => std_logic_vector'(x"00000000"),
  6023 => std_logic_vector'(x"00000000"),
  6024 => std_logic_vector'(x"00000000"),
  6025 => std_logic_vector'(x"00000000"),
  6026 => std_logic_vector'(x"00000000"),
  6027 => std_logic_vector'(x"00000000"),
  6028 => std_logic_vector'(x"00000000"),
  6029 => std_logic_vector'(x"00000000"),
  6030 => std_logic_vector'(x"00000000"),
  6031 => std_logic_vector'(x"00000000"),
  6032 => std_logic_vector'(x"00000000"),
  6033 => std_logic_vector'(x"00000000"),
  6034 => std_logic_vector'(x"00000000"),
  6035 => std_logic_vector'(x"00000000"),
  6036 => std_logic_vector'(x"00000000"),
  6037 => std_logic_vector'(x"00000000"),
  6038 => std_logic_vector'(x"00000000"),
  6039 => std_logic_vector'(x"00000000"),
  6040 => std_logic_vector'(x"00000000"),
  6041 => std_logic_vector'(x"00000000"),
  6042 => std_logic_vector'(x"00000000"),
  6043 => std_logic_vector'(x"00000000"),
  6044 => std_logic_vector'(x"00000000"),
  6045 => std_logic_vector'(x"00000000"),
  6046 => std_logic_vector'(x"00000000"),
  6047 => std_logic_vector'(x"00000000"),
  6048 => std_logic_vector'(x"00000000"),
  6049 => std_logic_vector'(x"00000000"),
  6050 => std_logic_vector'(x"00000000"),
  6051 => std_logic_vector'(x"00000000"),
  6052 => std_logic_vector'(x"00000000"),
  6053 => std_logic_vector'(x"00000000"),
  6054 => std_logic_vector'(x"00000000"),
  6055 => std_logic_vector'(x"00000000"),
  6056 => std_logic_vector'(x"00000000"),
  6057 => std_logic_vector'(x"00000000"),
  6058 => std_logic_vector'(x"00000000"),
  6059 => std_logic_vector'(x"00000000"),
  6060 => std_logic_vector'(x"00000000"),
  6061 => std_logic_vector'(x"00000000"),
  6062 => std_logic_vector'(x"00000000"),
  6063 => std_logic_vector'(x"00000000"),
  6064 => std_logic_vector'(x"00000000"),
  6065 => std_logic_vector'(x"00000000"),
  6066 => std_logic_vector'(x"00000000"),
  6067 => std_logic_vector'(x"00000000"),
  6068 => std_logic_vector'(x"00000000"),
  6069 => std_logic_vector'(x"00000000"),
  6070 => std_logic_vector'(x"00000000"),
  6071 => std_logic_vector'(x"00000000"),
  6072 => std_logic_vector'(x"00000000"),
  6073 => std_logic_vector'(x"00000000"),
  6074 => std_logic_vector'(x"00000000"),
  6075 => std_logic_vector'(x"00000000"),
  6076 => std_logic_vector'(x"00000000"),
  6077 => std_logic_vector'(x"00000000"),
  6078 => std_logic_vector'(x"00000000"),
  6079 => std_logic_vector'(x"00000000"),
  6080 => std_logic_vector'(x"00000000"),
  6081 => std_logic_vector'(x"00000000"),
  6082 => std_logic_vector'(x"00000000"),
  6083 => std_logic_vector'(x"00000000"),
  6084 => std_logic_vector'(x"00000000"),
  6085 => std_logic_vector'(x"00000000"),
  6086 => std_logic_vector'(x"00000000"),
  6087 => std_logic_vector'(x"00000000"),
  6088 => std_logic_vector'(x"00000000"),
  6089 => std_logic_vector'(x"00000000"),
  6090 => std_logic_vector'(x"00000000"),
  6091 => std_logic_vector'(x"00000000"),
  6092 => std_logic_vector'(x"00000000"),
  6093 => std_logic_vector'(x"00000000"),
  6094 => std_logic_vector'(x"00000000"),
  6095 => std_logic_vector'(x"00000000"),
  6096 => std_logic_vector'(x"00000000"),
  6097 => std_logic_vector'(x"00000000"),
  6098 => std_logic_vector'(x"00000000"),
  6099 => std_logic_vector'(x"00000000"),
  6100 => std_logic_vector'(x"00000000"),
  6101 => std_logic_vector'(x"00000000"),
  6102 => std_logic_vector'(x"00000000"),
  6103 => std_logic_vector'(x"00000000"),
  6104 => std_logic_vector'(x"00000000"),
  6105 => std_logic_vector'(x"00000000"),
  6106 => std_logic_vector'(x"00000000"),
  6107 => std_logic_vector'(x"00000000"),
  6108 => std_logic_vector'(x"00000000"),
  6109 => std_logic_vector'(x"00000000"),
  6110 => std_logic_vector'(x"00000000"),
  6111 => std_logic_vector'(x"00000000"),
  6112 => std_logic_vector'(x"00000000"),
  6113 => std_logic_vector'(x"00000000"),
  6114 => std_logic_vector'(x"00000000"),
  6115 => std_logic_vector'(x"00000000"),
  6116 => std_logic_vector'(x"00000000"),
  6117 => std_logic_vector'(x"00000000"),
  6118 => std_logic_vector'(x"00000000"),
  6119 => std_logic_vector'(x"00000000"),
  6120 => std_logic_vector'(x"00000000"),
  6121 => std_logic_vector'(x"00000000"),
  6122 => std_logic_vector'(x"00000000"),
  6123 => std_logic_vector'(x"00000000"),
  6124 => std_logic_vector'(x"00000000"),
  6125 => std_logic_vector'(x"00000000"),
  6126 => std_logic_vector'(x"00000000"),
  6127 => std_logic_vector'(x"00000000"),
  6128 => std_logic_vector'(x"00000000"),
  6129 => std_logic_vector'(x"00000000"),
  6130 => std_logic_vector'(x"00000000"),
  6131 => std_logic_vector'(x"00000000"),
  6132 => std_logic_vector'(x"00000000"),
  6133 => std_logic_vector'(x"00000000"),
  6134 => std_logic_vector'(x"00000000"),
  6135 => std_logic_vector'(x"00000000"),
  6136 => std_logic_vector'(x"00000000"),
  6137 => std_logic_vector'(x"00000000"),
  6138 => std_logic_vector'(x"00000000"),
  6139 => std_logic_vector'(x"00000000"),
  6140 => std_logic_vector'(x"00000000"),
  6141 => std_logic_vector'(x"00000000"),
  6142 => std_logic_vector'(x"00000000"),
  6143 => std_logic_vector'(x"00000000"),
  6144 => std_logic_vector'(x"00000000"),
  6145 => std_logic_vector'(x"00000000"),
  6146 => std_logic_vector'(x"00000000"),
  6147 => std_logic_vector'(x"00000000"),
  6148 => std_logic_vector'(x"00000000"),
  6149 => std_logic_vector'(x"00000000"),
  6150 => std_logic_vector'(x"00000000"),
  6151 => std_logic_vector'(x"00000000"),
  6152 => std_logic_vector'(x"00000000"),
  6153 => std_logic_vector'(x"00000000"),
  6154 => std_logic_vector'(x"00000000"),
  6155 => std_logic_vector'(x"00000000"),
  6156 => std_logic_vector'(x"00000000"),
  6157 => std_logic_vector'(x"00000000"),
  6158 => std_logic_vector'(x"00000000"),
  6159 => std_logic_vector'(x"00000000"),
  6160 => std_logic_vector'(x"00000000"),
  6161 => std_logic_vector'(x"00000000"),
  6162 => std_logic_vector'(x"00000000"),
  6163 => std_logic_vector'(x"00000000"),
  6164 => std_logic_vector'(x"00000000"),
  6165 => std_logic_vector'(x"00000000"),
  6166 => std_logic_vector'(x"00000000"),
  6167 => std_logic_vector'(x"00000000"),
  6168 => std_logic_vector'(x"00000000"),
  6169 => std_logic_vector'(x"00000000"),
  6170 => std_logic_vector'(x"00000000"),
  6171 => std_logic_vector'(x"00000000"),
  6172 => std_logic_vector'(x"00000000"),
  6173 => std_logic_vector'(x"00000000"),
  6174 => std_logic_vector'(x"00000000"),
  6175 => std_logic_vector'(x"00000000"),
  6176 => std_logic_vector'(x"00000000"),
  6177 => std_logic_vector'(x"00000000"),
  6178 => std_logic_vector'(x"00000000"),
  6179 => std_logic_vector'(x"00000000"),
  6180 => std_logic_vector'(x"00000000"),
  6181 => std_logic_vector'(x"00000000"),
  6182 => std_logic_vector'(x"00000000"),
  6183 => std_logic_vector'(x"00000000"),
  6184 => std_logic_vector'(x"00000000"),
  6185 => std_logic_vector'(x"00000000"),
  6186 => std_logic_vector'(x"00000000"),
  6187 => std_logic_vector'(x"00000000"),
  6188 => std_logic_vector'(x"00000000"),
  6189 => std_logic_vector'(x"00000000"),
  6190 => std_logic_vector'(x"00000000"),
  6191 => std_logic_vector'(x"00000000"),
  6192 => std_logic_vector'(x"00000000"),
  6193 => std_logic_vector'(x"00000000"),
  6194 => std_logic_vector'(x"00000000"),
  6195 => std_logic_vector'(x"00000000"),
  6196 => std_logic_vector'(x"00000000"),
  6197 => std_logic_vector'(x"00000000"),
  6198 => std_logic_vector'(x"00000000"),
  6199 => std_logic_vector'(x"00000000"),
  6200 => std_logic_vector'(x"00000000"),
  6201 => std_logic_vector'(x"00000000"),
  6202 => std_logic_vector'(x"00000000"),
  6203 => std_logic_vector'(x"00000000"),
  6204 => std_logic_vector'(x"00000000"),
  6205 => std_logic_vector'(x"00000000"),
  6206 => std_logic_vector'(x"00000000"),
  6207 => std_logic_vector'(x"00000000"),
  6208 => std_logic_vector'(x"00000000"),
  6209 => std_logic_vector'(x"00000000"),
  6210 => std_logic_vector'(x"00000000"),
  6211 => std_logic_vector'(x"00000000"),
  6212 => std_logic_vector'(x"00000000"),
  6213 => std_logic_vector'(x"00000000"),
  6214 => std_logic_vector'(x"00000000"),
  6215 => std_logic_vector'(x"00000000"),
  6216 => std_logic_vector'(x"00000000"),
  6217 => std_logic_vector'(x"00000000"),
  6218 => std_logic_vector'(x"00000000"),
  6219 => std_logic_vector'(x"00000000"),
  6220 => std_logic_vector'(x"00000000"),
  6221 => std_logic_vector'(x"00000000"),
  6222 => std_logic_vector'(x"00000000"),
  6223 => std_logic_vector'(x"00000000"),
  6224 => std_logic_vector'(x"00000000"),
  6225 => std_logic_vector'(x"00000000"),
  6226 => std_logic_vector'(x"00000000"),
  6227 => std_logic_vector'(x"00000000"),
  6228 => std_logic_vector'(x"00000000"),
  6229 => std_logic_vector'(x"00000000"),
  6230 => std_logic_vector'(x"00000000"),
  6231 => std_logic_vector'(x"00000000"),
  6232 => std_logic_vector'(x"00000000"),
  6233 => std_logic_vector'(x"00000000"),
  6234 => std_logic_vector'(x"00000000"),
  6235 => std_logic_vector'(x"00000000"),
  6236 => std_logic_vector'(x"00000000"),
  6237 => std_logic_vector'(x"00000000"),
  6238 => std_logic_vector'(x"00000000"),
  6239 => std_logic_vector'(x"00000000"),
  6240 => std_logic_vector'(x"00000000"),
  6241 => std_logic_vector'(x"00000000"),
  6242 => std_logic_vector'(x"00000000"),
  6243 => std_logic_vector'(x"00000000"),
  6244 => std_logic_vector'(x"00000000"),
  6245 => std_logic_vector'(x"00000000"),
  6246 => std_logic_vector'(x"00000000"),
  6247 => std_logic_vector'(x"00000000"),
  6248 => std_logic_vector'(x"00000000"),
  6249 => std_logic_vector'(x"00000000"),
  6250 => std_logic_vector'(x"00000000"),
  6251 => std_logic_vector'(x"00000000"),
  6252 => std_logic_vector'(x"00000000"),
  6253 => std_logic_vector'(x"00000000"),
  6254 => std_logic_vector'(x"00000000"),
  6255 => std_logic_vector'(x"00000000"),
  6256 => std_logic_vector'(x"00000000"),
  6257 => std_logic_vector'(x"00000000"),
  6258 => std_logic_vector'(x"00000000"),
  6259 => std_logic_vector'(x"00000000"),
  6260 => std_logic_vector'(x"00000000"),
  6261 => std_logic_vector'(x"00000000"),
  6262 => std_logic_vector'(x"00000000"),
  6263 => std_logic_vector'(x"00000000"),
  6264 => std_logic_vector'(x"00000000"),
  6265 => std_logic_vector'(x"00000000"),
  6266 => std_logic_vector'(x"00000000"),
  6267 => std_logic_vector'(x"00000000"),
  6268 => std_logic_vector'(x"00000000"),
  6269 => std_logic_vector'(x"00000000"),
  6270 => std_logic_vector'(x"00000000"),
  6271 => std_logic_vector'(x"00000000"),
  6272 => std_logic_vector'(x"00000000"),
  6273 => std_logic_vector'(x"00000000"),
  6274 => std_logic_vector'(x"00000000"),
  6275 => std_logic_vector'(x"00000000"),
  6276 => std_logic_vector'(x"00000000"),
  6277 => std_logic_vector'(x"00000000"),
  6278 => std_logic_vector'(x"00000000"),
  6279 => std_logic_vector'(x"00000000"),
  6280 => std_logic_vector'(x"00000000"),
  6281 => std_logic_vector'(x"00000000"),
  6282 => std_logic_vector'(x"00000000"),
  6283 => std_logic_vector'(x"00000000"),
  6284 => std_logic_vector'(x"00000000"),
  6285 => std_logic_vector'(x"00000000"),
  6286 => std_logic_vector'(x"00000000"),
  6287 => std_logic_vector'(x"00000000"),
  6288 => std_logic_vector'(x"00000000"),
  6289 => std_logic_vector'(x"00000000"),
  6290 => std_logic_vector'(x"00000000"),
  6291 => std_logic_vector'(x"00000000"),
  6292 => std_logic_vector'(x"00000000"),
  6293 => std_logic_vector'(x"00000000"),
  6294 => std_logic_vector'(x"00000000"),
  6295 => std_logic_vector'(x"00000000"),
  6296 => std_logic_vector'(x"00000000"),
  6297 => std_logic_vector'(x"00000000"),
  6298 => std_logic_vector'(x"00000000"),
  6299 => std_logic_vector'(x"00000000"),
  6300 => std_logic_vector'(x"00000000"),
  6301 => std_logic_vector'(x"00000000"),
  6302 => std_logic_vector'(x"00000000"),
  6303 => std_logic_vector'(x"00000000"),
  6304 => std_logic_vector'(x"00000000"),
  6305 => std_logic_vector'(x"00000000"),
  6306 => std_logic_vector'(x"00000000"),
  6307 => std_logic_vector'(x"00000000"),
  6308 => std_logic_vector'(x"00000000"),
  6309 => std_logic_vector'(x"00000000"),
  6310 => std_logic_vector'(x"00000000"),
  6311 => std_logic_vector'(x"00000000"),
  6312 => std_logic_vector'(x"00000000"),
  6313 => std_logic_vector'(x"00000000"),
  6314 => std_logic_vector'(x"00000000"),
  6315 => std_logic_vector'(x"00000000"),
  6316 => std_logic_vector'(x"00000000"),
  6317 => std_logic_vector'(x"00000000"),
  6318 => std_logic_vector'(x"00000000"),
  6319 => std_logic_vector'(x"00000000"),
  6320 => std_logic_vector'(x"00000000"),
  6321 => std_logic_vector'(x"00000000"),
  6322 => std_logic_vector'(x"00000000"),
  6323 => std_logic_vector'(x"00000000"),
  6324 => std_logic_vector'(x"00000000"),
  6325 => std_logic_vector'(x"00000000"),
  6326 => std_logic_vector'(x"00000000"),
  6327 => std_logic_vector'(x"00000000"),
  6328 => std_logic_vector'(x"00000000"),
  6329 => std_logic_vector'(x"00000000"),
  6330 => std_logic_vector'(x"00000000"),
  6331 => std_logic_vector'(x"00000000"),
  6332 => std_logic_vector'(x"00000000"),
  6333 => std_logic_vector'(x"00000000"),
  6334 => std_logic_vector'(x"00000000"),
  6335 => std_logic_vector'(x"00000000"),
  6336 => std_logic_vector'(x"00000000"),
  6337 => std_logic_vector'(x"00000000"),
  6338 => std_logic_vector'(x"00000000"),
  6339 => std_logic_vector'(x"00000000"),
  6340 => std_logic_vector'(x"00000000"),
  6341 => std_logic_vector'(x"00000000"),
  6342 => std_logic_vector'(x"00000000"),
  6343 => std_logic_vector'(x"00000000"),
  6344 => std_logic_vector'(x"00000000"),
  6345 => std_logic_vector'(x"00000000"),
  6346 => std_logic_vector'(x"00000000"),
  6347 => std_logic_vector'(x"00000000"),
  6348 => std_logic_vector'(x"00000000"),
  6349 => std_logic_vector'(x"00000000"),
  6350 => std_logic_vector'(x"00000000"),
  6351 => std_logic_vector'(x"00000000"),
  6352 => std_logic_vector'(x"00000000"),
  6353 => std_logic_vector'(x"00000000"),
  6354 => std_logic_vector'(x"00000000"),
  6355 => std_logic_vector'(x"00000000"),
  6356 => std_logic_vector'(x"00000000"),
  6357 => std_logic_vector'(x"00000000"),
  6358 => std_logic_vector'(x"00000000"),
  6359 => std_logic_vector'(x"00000000"),
  6360 => std_logic_vector'(x"00000000"),
  6361 => std_logic_vector'(x"00000000"),
  6362 => std_logic_vector'(x"00000000"),
  6363 => std_logic_vector'(x"00000000"),
  6364 => std_logic_vector'(x"00000000"),
  6365 => std_logic_vector'(x"00000000"),
  6366 => std_logic_vector'(x"00000000"),
  6367 => std_logic_vector'(x"00000000"),
  6368 => std_logic_vector'(x"00000000"),
  6369 => std_logic_vector'(x"00000000"),
  6370 => std_logic_vector'(x"00000000"),
  6371 => std_logic_vector'(x"00000000"),
  6372 => std_logic_vector'(x"00000000"),
  6373 => std_logic_vector'(x"00000000"),
  6374 => std_logic_vector'(x"00000000"),
  6375 => std_logic_vector'(x"00000000"),
  6376 => std_logic_vector'(x"00000000"),
  6377 => std_logic_vector'(x"00000000"),
  6378 => std_logic_vector'(x"00000000"),
  6379 => std_logic_vector'(x"00000000"),
  6380 => std_logic_vector'(x"00000000"),
  6381 => std_logic_vector'(x"00000000"),
  6382 => std_logic_vector'(x"00000000"),
  6383 => std_logic_vector'(x"00000000"),
  6384 => std_logic_vector'(x"00000000"),
  6385 => std_logic_vector'(x"00000000"),
  6386 => std_logic_vector'(x"00000000"),
  6387 => std_logic_vector'(x"00000000"),
  6388 => std_logic_vector'(x"00000000"),
  6389 => std_logic_vector'(x"00000000"),
  6390 => std_logic_vector'(x"00000000"),
  6391 => std_logic_vector'(x"00000000"),
  6392 => std_logic_vector'(x"00000000"),
  6393 => std_logic_vector'(x"00000000"),
  6394 => std_logic_vector'(x"00000000"),
  6395 => std_logic_vector'(x"00000000"),
  6396 => std_logic_vector'(x"00000000"),
  6397 => std_logic_vector'(x"00000000"),
  6398 => std_logic_vector'(x"00000000"),
  6399 => std_logic_vector'(x"00000000"),
  6400 => std_logic_vector'(x"00000000"),
  6401 => std_logic_vector'(x"00000000"),
  6402 => std_logic_vector'(x"00000000"),
  6403 => std_logic_vector'(x"00000000"),
  6404 => std_logic_vector'(x"00000000"),
  6405 => std_logic_vector'(x"00000000"),
  6406 => std_logic_vector'(x"00000000"),
  6407 => std_logic_vector'(x"00000000"),
  6408 => std_logic_vector'(x"00000000"),
  6409 => std_logic_vector'(x"00000000"),
  6410 => std_logic_vector'(x"00000000"),
  6411 => std_logic_vector'(x"00000000"),
  6412 => std_logic_vector'(x"00000000"),
  6413 => std_logic_vector'(x"00000000"),
  6414 => std_logic_vector'(x"00000000"),
  6415 => std_logic_vector'(x"00000000"),
  6416 => std_logic_vector'(x"00000000"),
  6417 => std_logic_vector'(x"00000000"),
  6418 => std_logic_vector'(x"00000000"),
  6419 => std_logic_vector'(x"00000000"),
  6420 => std_logic_vector'(x"00000000"),
  6421 => std_logic_vector'(x"00000000"),
  6422 => std_logic_vector'(x"00000000"),
  6423 => std_logic_vector'(x"00000000"),
  6424 => std_logic_vector'(x"00000000"),
  6425 => std_logic_vector'(x"00000000"),
  6426 => std_logic_vector'(x"00000000"),
  6427 => std_logic_vector'(x"00000000"),
  6428 => std_logic_vector'(x"00000000"),
  6429 => std_logic_vector'(x"00000000"),
  6430 => std_logic_vector'(x"00000000"),
  6431 => std_logic_vector'(x"00000000"),
  6432 => std_logic_vector'(x"00000000"),
  6433 => std_logic_vector'(x"00000000"),
  6434 => std_logic_vector'(x"00000000"),
  6435 => std_logic_vector'(x"00000000"),
  6436 => std_logic_vector'(x"00000000"),
  6437 => std_logic_vector'(x"00000000"),
  6438 => std_logic_vector'(x"00000000"),
  6439 => std_logic_vector'(x"00000000"),
  6440 => std_logic_vector'(x"00000000"),
  6441 => std_logic_vector'(x"00000000"),
  6442 => std_logic_vector'(x"00000000"),
  6443 => std_logic_vector'(x"00000000"),
  6444 => std_logic_vector'(x"00000000"),
  6445 => std_logic_vector'(x"00000000"),
  6446 => std_logic_vector'(x"00000000"),
  6447 => std_logic_vector'(x"00000000"),
  6448 => std_logic_vector'(x"00000000"),
  6449 => std_logic_vector'(x"00000000"),
  6450 => std_logic_vector'(x"00000000"),
  6451 => std_logic_vector'(x"00000000"),
  6452 => std_logic_vector'(x"00000000"),
  6453 => std_logic_vector'(x"00000000"),
  6454 => std_logic_vector'(x"00000000"),
  6455 => std_logic_vector'(x"00000000"),
  6456 => std_logic_vector'(x"00000000"),
  6457 => std_logic_vector'(x"00000000"),
  6458 => std_logic_vector'(x"00000000"),
  6459 => std_logic_vector'(x"00000000"),
  6460 => std_logic_vector'(x"00000000"),
  6461 => std_logic_vector'(x"00000000"),
  6462 => std_logic_vector'(x"00000000"),
  6463 => std_logic_vector'(x"00000000"),
  6464 => std_logic_vector'(x"00000000"),
  6465 => std_logic_vector'(x"00000000"),
  6466 => std_logic_vector'(x"00000000"),
  6467 => std_logic_vector'(x"00000000"),
  6468 => std_logic_vector'(x"00000000"),
  6469 => std_logic_vector'(x"00000000"),
  6470 => std_logic_vector'(x"00000000"),
  6471 => std_logic_vector'(x"00000000"),
  6472 => std_logic_vector'(x"00000000"),
  6473 => std_logic_vector'(x"00000000"),
  6474 => std_logic_vector'(x"00000000"),
  6475 => std_logic_vector'(x"00000000"),
  6476 => std_logic_vector'(x"00000000"),
  6477 => std_logic_vector'(x"00000000"),
  6478 => std_logic_vector'(x"00000000"),
  6479 => std_logic_vector'(x"00000000"),
  6480 => std_logic_vector'(x"00000000"),
  6481 => std_logic_vector'(x"00000000"),
  6482 => std_logic_vector'(x"00000000"),
  6483 => std_logic_vector'(x"00000000"),
  6484 => std_logic_vector'(x"00000000"),
  6485 => std_logic_vector'(x"00000000"),
  6486 => std_logic_vector'(x"00000000"),
  6487 => std_logic_vector'(x"00000000"),
  6488 => std_logic_vector'(x"00000000"),
  6489 => std_logic_vector'(x"00000000"),
  6490 => std_logic_vector'(x"00000000"),
  6491 => std_logic_vector'(x"00000000"),
  6492 => std_logic_vector'(x"00000000"),
  6493 => std_logic_vector'(x"00000000"),
  6494 => std_logic_vector'(x"00000000"),
  6495 => std_logic_vector'(x"00000000"),
  6496 => std_logic_vector'(x"00000000"),
  6497 => std_logic_vector'(x"00000000"),
  6498 => std_logic_vector'(x"00000000"),
  6499 => std_logic_vector'(x"00000000"),
  6500 => std_logic_vector'(x"00000000"),
  6501 => std_logic_vector'(x"00000000"),
  6502 => std_logic_vector'(x"00000000"),
  6503 => std_logic_vector'(x"00000000"),
  6504 => std_logic_vector'(x"00000000"),
  6505 => std_logic_vector'(x"00000000"),
  6506 => std_logic_vector'(x"00000000"),
  6507 => std_logic_vector'(x"00000000"),
  6508 => std_logic_vector'(x"00000000"),
  6509 => std_logic_vector'(x"00000000"),
  6510 => std_logic_vector'(x"00000000"),
  6511 => std_logic_vector'(x"00000000"),
  6512 => std_logic_vector'(x"00000000"),
  6513 => std_logic_vector'(x"00000000"),
  6514 => std_logic_vector'(x"00000000"),
  6515 => std_logic_vector'(x"00000000"),
  6516 => std_logic_vector'(x"00000000"),
  6517 => std_logic_vector'(x"00000000"),
  6518 => std_logic_vector'(x"00000000"),
  6519 => std_logic_vector'(x"00000000"),
  6520 => std_logic_vector'(x"00000000"),
  6521 => std_logic_vector'(x"00000000"),
  6522 => std_logic_vector'(x"00000000"),
  6523 => std_logic_vector'(x"00000000"),
  6524 => std_logic_vector'(x"00000000"),
  6525 => std_logic_vector'(x"00000000"),
  6526 => std_logic_vector'(x"00000000"),
  6527 => std_logic_vector'(x"00000000"),
  6528 => std_logic_vector'(x"00000000"),
  6529 => std_logic_vector'(x"00000000"),
  6530 => std_logic_vector'(x"00000000"),
  6531 => std_logic_vector'(x"00000000"),
  6532 => std_logic_vector'(x"00000000"),
  6533 => std_logic_vector'(x"00000000"),
  6534 => std_logic_vector'(x"00000000"),
  6535 => std_logic_vector'(x"00000000"),
  6536 => std_logic_vector'(x"00000000"),
  6537 => std_logic_vector'(x"00000000"),
  6538 => std_logic_vector'(x"00000000"),
  6539 => std_logic_vector'(x"00000000"),
  6540 => std_logic_vector'(x"00000000"),
  6541 => std_logic_vector'(x"00000000"),
  6542 => std_logic_vector'(x"00000000"),
  6543 => std_logic_vector'(x"00000000"),
  6544 => std_logic_vector'(x"00000000"),
  6545 => std_logic_vector'(x"00000000"),
  6546 => std_logic_vector'(x"00000000"),
  6547 => std_logic_vector'(x"00000000"),
  6548 => std_logic_vector'(x"00000000"),
  6549 => std_logic_vector'(x"00000000"),
  6550 => std_logic_vector'(x"00000000"),
  6551 => std_logic_vector'(x"00000000"),
  6552 => std_logic_vector'(x"00000000"),
  6553 => std_logic_vector'(x"00000000"),
  6554 => std_logic_vector'(x"00000000"),
  6555 => std_logic_vector'(x"00000000"),
  6556 => std_logic_vector'(x"00000000"),
  6557 => std_logic_vector'(x"00000000"),
  6558 => std_logic_vector'(x"00000000"),
  6559 => std_logic_vector'(x"00000000"),
  6560 => std_logic_vector'(x"00000000"),
  6561 => std_logic_vector'(x"00000000"),
  6562 => std_logic_vector'(x"00000000"),
  6563 => std_logic_vector'(x"00000000"),
  6564 => std_logic_vector'(x"00000000"),
  6565 => std_logic_vector'(x"00000000"),
  6566 => std_logic_vector'(x"00000000"),
  6567 => std_logic_vector'(x"00000000"),
  6568 => std_logic_vector'(x"00000000"),
  6569 => std_logic_vector'(x"00000000"),
  6570 => std_logic_vector'(x"00000000"),
  6571 => std_logic_vector'(x"00000000"),
  6572 => std_logic_vector'(x"00000000"),
  6573 => std_logic_vector'(x"00000000"),
  6574 => std_logic_vector'(x"00000000"),
  6575 => std_logic_vector'(x"00000000"),
  6576 => std_logic_vector'(x"00000000"),
  6577 => std_logic_vector'(x"00000000"),
  6578 => std_logic_vector'(x"00000000"),
  6579 => std_logic_vector'(x"00000000"),
  6580 => std_logic_vector'(x"00000000"),
  6581 => std_logic_vector'(x"00000000"),
  6582 => std_logic_vector'(x"00000000"),
  6583 => std_logic_vector'(x"00000000"),
  6584 => std_logic_vector'(x"00000000"),
  6585 => std_logic_vector'(x"00000000"),
  6586 => std_logic_vector'(x"00000000"),
  6587 => std_logic_vector'(x"00000000"),
  6588 => std_logic_vector'(x"00000000"),
  6589 => std_logic_vector'(x"00000000"),
  6590 => std_logic_vector'(x"00000000"),
  6591 => std_logic_vector'(x"00000000"),
  6592 => std_logic_vector'(x"00000000"),
  6593 => std_logic_vector'(x"00000000"),
  6594 => std_logic_vector'(x"00000000"),
  6595 => std_logic_vector'(x"00000000"),
  6596 => std_logic_vector'(x"00000000"),
  6597 => std_logic_vector'(x"00000000"),
  6598 => std_logic_vector'(x"00000000"),
  6599 => std_logic_vector'(x"00000000"),
  6600 => std_logic_vector'(x"00000000"),
  6601 => std_logic_vector'(x"00000000"),
  6602 => std_logic_vector'(x"00000000"),
  6603 => std_logic_vector'(x"00000000"),
  6604 => std_logic_vector'(x"00000000"),
  6605 => std_logic_vector'(x"00000000"),
  6606 => std_logic_vector'(x"00000000"),
  6607 => std_logic_vector'(x"00000000"),
  6608 => std_logic_vector'(x"00000000"),
  6609 => std_logic_vector'(x"00000000"),
  6610 => std_logic_vector'(x"00000000"),
  6611 => std_logic_vector'(x"00000000"),
  6612 => std_logic_vector'(x"00000000"),
  6613 => std_logic_vector'(x"00000000"),
  6614 => std_logic_vector'(x"00000000"),
  6615 => std_logic_vector'(x"00000000"),
  6616 => std_logic_vector'(x"00000000"),
  6617 => std_logic_vector'(x"00000000"),
  6618 => std_logic_vector'(x"00000000"),
  6619 => std_logic_vector'(x"00000000"),
  6620 => std_logic_vector'(x"00000000"),
  6621 => std_logic_vector'(x"00000000"),
  6622 => std_logic_vector'(x"00000000"),
  6623 => std_logic_vector'(x"00000000"),
  6624 => std_logic_vector'(x"00000000"),
  6625 => std_logic_vector'(x"00000000"),
  6626 => std_logic_vector'(x"00000000"),
  6627 => std_logic_vector'(x"00000000"),
  6628 => std_logic_vector'(x"00000000"),
  6629 => std_logic_vector'(x"00000000"),
  6630 => std_logic_vector'(x"00000000"),
  6631 => std_logic_vector'(x"00000000"),
  6632 => std_logic_vector'(x"00000000"),
  6633 => std_logic_vector'(x"00000000"),
  6634 => std_logic_vector'(x"00000000"),
  6635 => std_logic_vector'(x"00000000"),
  6636 => std_logic_vector'(x"00000000"),
  6637 => std_logic_vector'(x"00000000"),
  6638 => std_logic_vector'(x"00000000"),
  6639 => std_logic_vector'(x"00000000"),
  6640 => std_logic_vector'(x"00000000"),
  6641 => std_logic_vector'(x"00000000"),
  6642 => std_logic_vector'(x"00000000"),
  6643 => std_logic_vector'(x"00000000"),
  6644 => std_logic_vector'(x"00000000"),
  6645 => std_logic_vector'(x"00000000"),
  6646 => std_logic_vector'(x"00000000"),
  6647 => std_logic_vector'(x"00000000"),
  6648 => std_logic_vector'(x"00000000"),
  6649 => std_logic_vector'(x"00000000"),
  6650 => std_logic_vector'(x"00000000"),
  6651 => std_logic_vector'(x"00000000"),
  6652 => std_logic_vector'(x"00000000"),
  6653 => std_logic_vector'(x"00000000"),
  6654 => std_logic_vector'(x"00000000"),
  6655 => std_logic_vector'(x"00000000"),
  6656 => std_logic_vector'(x"00000000"),
  6657 => std_logic_vector'(x"00000000"),
  6658 => std_logic_vector'(x"00000000"),
  6659 => std_logic_vector'(x"00000000"),
  6660 => std_logic_vector'(x"00000000"),
  6661 => std_logic_vector'(x"00000000"),
  6662 => std_logic_vector'(x"00000000"),
  6663 => std_logic_vector'(x"00000000"),
  6664 => std_logic_vector'(x"00000000"),
  6665 => std_logic_vector'(x"00000000"),
  6666 => std_logic_vector'(x"00000000"),
  6667 => std_logic_vector'(x"00000000"),
  6668 => std_logic_vector'(x"00000000"),
  6669 => std_logic_vector'(x"00000000"),
  6670 => std_logic_vector'(x"00000000"),
  6671 => std_logic_vector'(x"00000000"),
  6672 => std_logic_vector'(x"00000000"),
  6673 => std_logic_vector'(x"00000000"),
  6674 => std_logic_vector'(x"00000000"),
  6675 => std_logic_vector'(x"00000000"),
  6676 => std_logic_vector'(x"00000000"),
  6677 => std_logic_vector'(x"00000000"),
  6678 => std_logic_vector'(x"00000000"),
  6679 => std_logic_vector'(x"00000000"),
  6680 => std_logic_vector'(x"00000000"),
  6681 => std_logic_vector'(x"00000000"),
  6682 => std_logic_vector'(x"00000000"),
  6683 => std_logic_vector'(x"00000000"),
  6684 => std_logic_vector'(x"00000000"),
  6685 => std_logic_vector'(x"00000000"),
  6686 => std_logic_vector'(x"00000000"),
  6687 => std_logic_vector'(x"00000000"),
  6688 => std_logic_vector'(x"00000000"),
  6689 => std_logic_vector'(x"00000000"),
  6690 => std_logic_vector'(x"00000000"),
  6691 => std_logic_vector'(x"00000000"),
  6692 => std_logic_vector'(x"00000000"),
  6693 => std_logic_vector'(x"00000000"),
  6694 => std_logic_vector'(x"00000000"),
  6695 => std_logic_vector'(x"00000000"),
  6696 => std_logic_vector'(x"00000000"),
  6697 => std_logic_vector'(x"00000000"),
  6698 => std_logic_vector'(x"00000000"),
  6699 => std_logic_vector'(x"00000000"),
  6700 => std_logic_vector'(x"00000000"),
  6701 => std_logic_vector'(x"00000000"),
  6702 => std_logic_vector'(x"00000000"),
  6703 => std_logic_vector'(x"00000000"),
  6704 => std_logic_vector'(x"00000000"),
  6705 => std_logic_vector'(x"00000000"),
  6706 => std_logic_vector'(x"00000000"),
  6707 => std_logic_vector'(x"00000000"),
  6708 => std_logic_vector'(x"00000000"),
  6709 => std_logic_vector'(x"00000000"),
  6710 => std_logic_vector'(x"00000000"),
  6711 => std_logic_vector'(x"00000000"),
  6712 => std_logic_vector'(x"00000000"),
  6713 => std_logic_vector'(x"00000000"),
  6714 => std_logic_vector'(x"00000000"),
  6715 => std_logic_vector'(x"00000000"),
  6716 => std_logic_vector'(x"00000000"),
  6717 => std_logic_vector'(x"00000000"),
  6718 => std_logic_vector'(x"00000000"),
  6719 => std_logic_vector'(x"00000000"),
  6720 => std_logic_vector'(x"00000000"),
  6721 => std_logic_vector'(x"00000000"),
  6722 => std_logic_vector'(x"00000000"),
  6723 => std_logic_vector'(x"00000000"),
  6724 => std_logic_vector'(x"00000000"),
  6725 => std_logic_vector'(x"00000000"),
  6726 => std_logic_vector'(x"00000000"),
  6727 => std_logic_vector'(x"00000000"),
  6728 => std_logic_vector'(x"00000000"),
  6729 => std_logic_vector'(x"00000000"),
  6730 => std_logic_vector'(x"00000000"),
  6731 => std_logic_vector'(x"00000000"),
  6732 => std_logic_vector'(x"00000000"),
  6733 => std_logic_vector'(x"00000000"),
  6734 => std_logic_vector'(x"00000000"),
  6735 => std_logic_vector'(x"00000000"),
  6736 => std_logic_vector'(x"00000000"),
  6737 => std_logic_vector'(x"00000000"),
  6738 => std_logic_vector'(x"00000000"),
  6739 => std_logic_vector'(x"00000000"),
  6740 => std_logic_vector'(x"00000000"),
  6741 => std_logic_vector'(x"00000000"),
  6742 => std_logic_vector'(x"00000000"),
  6743 => std_logic_vector'(x"00000000"),
  6744 => std_logic_vector'(x"00000000"),
  6745 => std_logic_vector'(x"00000000"),
  6746 => std_logic_vector'(x"00000000"),
  6747 => std_logic_vector'(x"00000000"),
  6748 => std_logic_vector'(x"00000000"),
  6749 => std_logic_vector'(x"00000000"),
  6750 => std_logic_vector'(x"00000000"),
  6751 => std_logic_vector'(x"00000000"),
  6752 => std_logic_vector'(x"00000000"),
  6753 => std_logic_vector'(x"00000000"),
  6754 => std_logic_vector'(x"00000000"),
  6755 => std_logic_vector'(x"00000000"),
  6756 => std_logic_vector'(x"00000000"),
  6757 => std_logic_vector'(x"00000000"),
  6758 => std_logic_vector'(x"00000000"),
  6759 => std_logic_vector'(x"00000000"),
  6760 => std_logic_vector'(x"00000000"),
  6761 => std_logic_vector'(x"00000000"),
  6762 => std_logic_vector'(x"00000000"),
  6763 => std_logic_vector'(x"00000000"),
  6764 => std_logic_vector'(x"00000000"),
  6765 => std_logic_vector'(x"00000000"),
  6766 => std_logic_vector'(x"00000000"),
  6767 => std_logic_vector'(x"00000000"),
  6768 => std_logic_vector'(x"00000000"),
  6769 => std_logic_vector'(x"00000000"),
  6770 => std_logic_vector'(x"00000000"),
  6771 => std_logic_vector'(x"00000000"),
  6772 => std_logic_vector'(x"00000000"),
  6773 => std_logic_vector'(x"00000000"),
  6774 => std_logic_vector'(x"00000000"),
  6775 => std_logic_vector'(x"00000000"),
  6776 => std_logic_vector'(x"00000000"),
  6777 => std_logic_vector'(x"00000000"),
  6778 => std_logic_vector'(x"00000000"),
  6779 => std_logic_vector'(x"00000000"),
  6780 => std_logic_vector'(x"00000000"),
  6781 => std_logic_vector'(x"00000000"),
  6782 => std_logic_vector'(x"00000000"),
  6783 => std_logic_vector'(x"00000000"),
  6784 => std_logic_vector'(x"00000000"),
  6785 => std_logic_vector'(x"00000000"),
  6786 => std_logic_vector'(x"00000000"),
  6787 => std_logic_vector'(x"00000000"),
  6788 => std_logic_vector'(x"00000000"),
  6789 => std_logic_vector'(x"00000000"),
  6790 => std_logic_vector'(x"00000000"),
  6791 => std_logic_vector'(x"00000000"),
  6792 => std_logic_vector'(x"00000000"),
  6793 => std_logic_vector'(x"00000000"),
  6794 => std_logic_vector'(x"00000000"),
  6795 => std_logic_vector'(x"00000000"),
  6796 => std_logic_vector'(x"00000000"),
  6797 => std_logic_vector'(x"00000000"),
  6798 => std_logic_vector'(x"00000000"),
  6799 => std_logic_vector'(x"00000000"),
  6800 => std_logic_vector'(x"00000000"),
  6801 => std_logic_vector'(x"00000000"),
  6802 => std_logic_vector'(x"00000000"),
  6803 => std_logic_vector'(x"00000000"),
  6804 => std_logic_vector'(x"00000000"),
  6805 => std_logic_vector'(x"00000000"),
  6806 => std_logic_vector'(x"00000000"),
  6807 => std_logic_vector'(x"00000000"),
  6808 => std_logic_vector'(x"00000000"),
  6809 => std_logic_vector'(x"00000000"),
  6810 => std_logic_vector'(x"00000000"),
  6811 => std_logic_vector'(x"00000000"),
  6812 => std_logic_vector'(x"00000000"),
  6813 => std_logic_vector'(x"00000000"),
  6814 => std_logic_vector'(x"00000000"),
  6815 => std_logic_vector'(x"00000000"),
  6816 => std_logic_vector'(x"00000000"),
  6817 => std_logic_vector'(x"00000000"),
  6818 => std_logic_vector'(x"00000000"),
  6819 => std_logic_vector'(x"00000000"),
  6820 => std_logic_vector'(x"00000000"),
  6821 => std_logic_vector'(x"00000000"),
  6822 => std_logic_vector'(x"00000000"),
  6823 => std_logic_vector'(x"00000000"),
  6824 => std_logic_vector'(x"00000000"),
  6825 => std_logic_vector'(x"00000000"),
  6826 => std_logic_vector'(x"00000000"),
  6827 => std_logic_vector'(x"00000000"),
  6828 => std_logic_vector'(x"00000000"),
  6829 => std_logic_vector'(x"00000000"),
  6830 => std_logic_vector'(x"00000000"),
  6831 => std_logic_vector'(x"00000000"),
  6832 => std_logic_vector'(x"00000000"),
  6833 => std_logic_vector'(x"00000000"),
  6834 => std_logic_vector'(x"00000000"),
  6835 => std_logic_vector'(x"00000000"),
  6836 => std_logic_vector'(x"00000000"),
  6837 => std_logic_vector'(x"00000000"),
  6838 => std_logic_vector'(x"00000000"),
  6839 => std_logic_vector'(x"00000000"),
  6840 => std_logic_vector'(x"00000000"),
  6841 => std_logic_vector'(x"00000000"),
  6842 => std_logic_vector'(x"00000000"),
  6843 => std_logic_vector'(x"00000000"),
  6844 => std_logic_vector'(x"00000000"),
  6845 => std_logic_vector'(x"00000000"),
  6846 => std_logic_vector'(x"00000000"),
  6847 => std_logic_vector'(x"00000000"),
  6848 => std_logic_vector'(x"00000000"),
  6849 => std_logic_vector'(x"00000000"),
  6850 => std_logic_vector'(x"00000000"),
  6851 => std_logic_vector'(x"00000000"),
  6852 => std_logic_vector'(x"00000000"),
  6853 => std_logic_vector'(x"00000000"),
  6854 => std_logic_vector'(x"00000000"),
  6855 => std_logic_vector'(x"00000000"),
  6856 => std_logic_vector'(x"00000000"),
  6857 => std_logic_vector'(x"00000000"),
  6858 => std_logic_vector'(x"00000000"),
  6859 => std_logic_vector'(x"00000000"),
  6860 => std_logic_vector'(x"00000000"),
  6861 => std_logic_vector'(x"00000000"),
  6862 => std_logic_vector'(x"00000000"),
  6863 => std_logic_vector'(x"00000000"),
  6864 => std_logic_vector'(x"00000000"),
  6865 => std_logic_vector'(x"00000000"),
  6866 => std_logic_vector'(x"00000000"),
  6867 => std_logic_vector'(x"00000000"),
  6868 => std_logic_vector'(x"00000000"),
  6869 => std_logic_vector'(x"00000000"),
  6870 => std_logic_vector'(x"00000000"),
  6871 => std_logic_vector'(x"00000000"),
  6872 => std_logic_vector'(x"00000000"),
  6873 => std_logic_vector'(x"00000000"),
  6874 => std_logic_vector'(x"00000000"),
  6875 => std_logic_vector'(x"00000000"),
  6876 => std_logic_vector'(x"00000000"),
  6877 => std_logic_vector'(x"00000000"),
  6878 => std_logic_vector'(x"00000000"),
  6879 => std_logic_vector'(x"00000000"),
  6880 => std_logic_vector'(x"00000000"),
  6881 => std_logic_vector'(x"00000000"),
  6882 => std_logic_vector'(x"00000000"),
  6883 => std_logic_vector'(x"00000000"),
  6884 => std_logic_vector'(x"00000000"),
  6885 => std_logic_vector'(x"00000000"),
  6886 => std_logic_vector'(x"00000000"),
  6887 => std_logic_vector'(x"00000000"),
  6888 => std_logic_vector'(x"00000000"),
  6889 => std_logic_vector'(x"00000000"),
  6890 => std_logic_vector'(x"00000000"),
  6891 => std_logic_vector'(x"00000000"),
  6892 => std_logic_vector'(x"00000000"),
  6893 => std_logic_vector'(x"00000000"),
  6894 => std_logic_vector'(x"00000000"),
  6895 => std_logic_vector'(x"00000000"),
  6896 => std_logic_vector'(x"00000000"),
  6897 => std_logic_vector'(x"00000000"),
  6898 => std_logic_vector'(x"00000000"),
  6899 => std_logic_vector'(x"00000000"),
  6900 => std_logic_vector'(x"00000000"),
  6901 => std_logic_vector'(x"00000000"),
  6902 => std_logic_vector'(x"00000000"),
  6903 => std_logic_vector'(x"00000000"),
  6904 => std_logic_vector'(x"00000000"),
  6905 => std_logic_vector'(x"00000000"),
  6906 => std_logic_vector'(x"00000000"),
  6907 => std_logic_vector'(x"00000000"),
  6908 => std_logic_vector'(x"00000000"),
  6909 => std_logic_vector'(x"00000000"),
  6910 => std_logic_vector'(x"00000000"),
  6911 => std_logic_vector'(x"00000000"),
  6912 => std_logic_vector'(x"00000000"),
  6913 => std_logic_vector'(x"00000000"),
  6914 => std_logic_vector'(x"00000000"),
  6915 => std_logic_vector'(x"00000000"),
  6916 => std_logic_vector'(x"00000000"),
  6917 => std_logic_vector'(x"00000000"),
  6918 => std_logic_vector'(x"00000000"),
  6919 => std_logic_vector'(x"00000000"),
  6920 => std_logic_vector'(x"00000000"),
  6921 => std_logic_vector'(x"00000000"),
  6922 => std_logic_vector'(x"00000000"),
  6923 => std_logic_vector'(x"00000000"),
  6924 => std_logic_vector'(x"00000000"),
  6925 => std_logic_vector'(x"00000000"),
  6926 => std_logic_vector'(x"00000000"),
  6927 => std_logic_vector'(x"00000000"),
  6928 => std_logic_vector'(x"00000000"),
  6929 => std_logic_vector'(x"00000000"),
  6930 => std_logic_vector'(x"00000000"),
  6931 => std_logic_vector'(x"00000000"),
  6932 => std_logic_vector'(x"00000000"),
  6933 => std_logic_vector'(x"00000000"),
  6934 => std_logic_vector'(x"00000000"),
  6935 => std_logic_vector'(x"00000000"),
  6936 => std_logic_vector'(x"00000000"),
  6937 => std_logic_vector'(x"00000000"),
  6938 => std_logic_vector'(x"00000000"),
  6939 => std_logic_vector'(x"00000000"),
  6940 => std_logic_vector'(x"00000000"),
  6941 => std_logic_vector'(x"00000000"),
  6942 => std_logic_vector'(x"00000000"),
  6943 => std_logic_vector'(x"00000000"),
  6944 => std_logic_vector'(x"00000000"),
  6945 => std_logic_vector'(x"00000000"),
  6946 => std_logic_vector'(x"00000000"),
  6947 => std_logic_vector'(x"00000000"),
  6948 => std_logic_vector'(x"00000000"),
  6949 => std_logic_vector'(x"00000000"),
  6950 => std_logic_vector'(x"00000000"),
  6951 => std_logic_vector'(x"00000000"),
  6952 => std_logic_vector'(x"00000000"),
  6953 => std_logic_vector'(x"00000000"),
  6954 => std_logic_vector'(x"00000000"),
  6955 => std_logic_vector'(x"00000000"),
  6956 => std_logic_vector'(x"00000000"),
  6957 => std_logic_vector'(x"00000000"),
  6958 => std_logic_vector'(x"00000000"),
  6959 => std_logic_vector'(x"00000000"),
  6960 => std_logic_vector'(x"00000000"),
  6961 => std_logic_vector'(x"00000000"),
  6962 => std_logic_vector'(x"00000000"),
  6963 => std_logic_vector'(x"00000000"),
  6964 => std_logic_vector'(x"00000000"),
  6965 => std_logic_vector'(x"00000000"),
  6966 => std_logic_vector'(x"00000000"),
  6967 => std_logic_vector'(x"00000000"),
  6968 => std_logic_vector'(x"00000000"),
  6969 => std_logic_vector'(x"00000000"),
  6970 => std_logic_vector'(x"00000000"),
  6971 => std_logic_vector'(x"00000000"),
  6972 => std_logic_vector'(x"00000000"),
  6973 => std_logic_vector'(x"00000000"),
  6974 => std_logic_vector'(x"00000000"),
  6975 => std_logic_vector'(x"00000000"),
  6976 => std_logic_vector'(x"00000000"),
  6977 => std_logic_vector'(x"00000000"),
  6978 => std_logic_vector'(x"00000000"),
  6979 => std_logic_vector'(x"00000000"),
  6980 => std_logic_vector'(x"00000000"),
  6981 => std_logic_vector'(x"00000000"),
  6982 => std_logic_vector'(x"00000000"),
  6983 => std_logic_vector'(x"00000000"),
  6984 => std_logic_vector'(x"00000000"),
  6985 => std_logic_vector'(x"00000000"),
  6986 => std_logic_vector'(x"00000000"),
  6987 => std_logic_vector'(x"00000000"),
  6988 => std_logic_vector'(x"00000000"),
  6989 => std_logic_vector'(x"00000000"),
  6990 => std_logic_vector'(x"00000000"),
  6991 => std_logic_vector'(x"00000000"),
  6992 => std_logic_vector'(x"00000000"),
  6993 => std_logic_vector'(x"00000000"),
  6994 => std_logic_vector'(x"00000000"),
  6995 => std_logic_vector'(x"00000000"),
  6996 => std_logic_vector'(x"00000000"),
  6997 => std_logic_vector'(x"00000000"),
  6998 => std_logic_vector'(x"00000000"),
  6999 => std_logic_vector'(x"00000000"),
  7000 => std_logic_vector'(x"00000000"),
  7001 => std_logic_vector'(x"00000000"),
  7002 => std_logic_vector'(x"00000000"),
  7003 => std_logic_vector'(x"00000000"),
  7004 => std_logic_vector'(x"00000000"),
  7005 => std_logic_vector'(x"00000000"),
  7006 => std_logic_vector'(x"00000000"),
  7007 => std_logic_vector'(x"00000000"),
  7008 => std_logic_vector'(x"00000000"),
  7009 => std_logic_vector'(x"00000000"),
  7010 => std_logic_vector'(x"00000000"),
  7011 => std_logic_vector'(x"00000000"),
  7012 => std_logic_vector'(x"00000000"),
  7013 => std_logic_vector'(x"00000000"),
  7014 => std_logic_vector'(x"00000000"),
  7015 => std_logic_vector'(x"00000000"),
  7016 => std_logic_vector'(x"00000000"),
  7017 => std_logic_vector'(x"00000000"),
  7018 => std_logic_vector'(x"00000000"),
  7019 => std_logic_vector'(x"00000000"),
  7020 => std_logic_vector'(x"00000000"),
  7021 => std_logic_vector'(x"00000000"),
  7022 => std_logic_vector'(x"00000000"),
  7023 => std_logic_vector'(x"00000000"),
  7024 => std_logic_vector'(x"00000000"),
  7025 => std_logic_vector'(x"00000000"),
  7026 => std_logic_vector'(x"00000000"),
  7027 => std_logic_vector'(x"00000000"),
  7028 => std_logic_vector'(x"00000000"),
  7029 => std_logic_vector'(x"00000000"),
  7030 => std_logic_vector'(x"00000000"),
  7031 => std_logic_vector'(x"00000000"),
  7032 => std_logic_vector'(x"00000000"),
  7033 => std_logic_vector'(x"00000000"),
  7034 => std_logic_vector'(x"00000000"),
  7035 => std_logic_vector'(x"00000000"),
  7036 => std_logic_vector'(x"00000000"),
  7037 => std_logic_vector'(x"00000000"),
  7038 => std_logic_vector'(x"00000000"),
  7039 => std_logic_vector'(x"00000000"),
  7040 => std_logic_vector'(x"00000000"),
  7041 => std_logic_vector'(x"00000000"),
  7042 => std_logic_vector'(x"00000000"),
  7043 => std_logic_vector'(x"00000000"),
  7044 => std_logic_vector'(x"00000000"),
  7045 => std_logic_vector'(x"00000000"),
  7046 => std_logic_vector'(x"00000000"),
  7047 => std_logic_vector'(x"00000000"),
  7048 => std_logic_vector'(x"00000000"),
  7049 => std_logic_vector'(x"00000000"),
  7050 => std_logic_vector'(x"00000000"),
  7051 => std_logic_vector'(x"00000000"),
  7052 => std_logic_vector'(x"00000000"),
  7053 => std_logic_vector'(x"00000000"),
  7054 => std_logic_vector'(x"00000000"),
  7055 => std_logic_vector'(x"00000000"),
  7056 => std_logic_vector'(x"00000000"),
  7057 => std_logic_vector'(x"00000000"),
  7058 => std_logic_vector'(x"00000000"),
  7059 => std_logic_vector'(x"00000000"),
  7060 => std_logic_vector'(x"00000000"),
  7061 => std_logic_vector'(x"00000000"),
  7062 => std_logic_vector'(x"00000000"),
  7063 => std_logic_vector'(x"00000000"),
  7064 => std_logic_vector'(x"00000000"),
  7065 => std_logic_vector'(x"00000000"),
  7066 => std_logic_vector'(x"00000000"),
  7067 => std_logic_vector'(x"00000000"),
  7068 => std_logic_vector'(x"00000000"),
  7069 => std_logic_vector'(x"00000000"),
  7070 => std_logic_vector'(x"00000000"),
  7071 => std_logic_vector'(x"00000000"),
  7072 => std_logic_vector'(x"00000000"),
  7073 => std_logic_vector'(x"00000000"),
  7074 => std_logic_vector'(x"00000000"),
  7075 => std_logic_vector'(x"00000000"),
  7076 => std_logic_vector'(x"00000000"),
  7077 => std_logic_vector'(x"00000000"),
  7078 => std_logic_vector'(x"00000000"),
  7079 => std_logic_vector'(x"00000000"),
  7080 => std_logic_vector'(x"00000000"),
  7081 => std_logic_vector'(x"00000000"),
  7082 => std_logic_vector'(x"00000000"),
  7083 => std_logic_vector'(x"00000000"),
  7084 => std_logic_vector'(x"00000000"),
  7085 => std_logic_vector'(x"00000000"),
  7086 => std_logic_vector'(x"00000000"),
  7087 => std_logic_vector'(x"00000000"),
  7088 => std_logic_vector'(x"00000000"),
  7089 => std_logic_vector'(x"00000000"),
  7090 => std_logic_vector'(x"00000000"),
  7091 => std_logic_vector'(x"00000000"),
  7092 => std_logic_vector'(x"00000000"),
  7093 => std_logic_vector'(x"00000000"),
  7094 => std_logic_vector'(x"00000000"),
  7095 => std_logic_vector'(x"00000000"),
  7096 => std_logic_vector'(x"00000000"),
  7097 => std_logic_vector'(x"00000000"),
  7098 => std_logic_vector'(x"00000000"),
  7099 => std_logic_vector'(x"00000000"),
  7100 => std_logic_vector'(x"00000000"),
  7101 => std_logic_vector'(x"00000000"),
  7102 => std_logic_vector'(x"00000000"),
  7103 => std_logic_vector'(x"00000000"),
  7104 => std_logic_vector'(x"00000000"),
  7105 => std_logic_vector'(x"00000000"),
  7106 => std_logic_vector'(x"00000000"),
  7107 => std_logic_vector'(x"00000000"),
  7108 => std_logic_vector'(x"00000000"),
  7109 => std_logic_vector'(x"00000000"),
  7110 => std_logic_vector'(x"00000000"),
  7111 => std_logic_vector'(x"00000000"),
  7112 => std_logic_vector'(x"00000000"),
  7113 => std_logic_vector'(x"00000000"),
  7114 => std_logic_vector'(x"00000000"),
  7115 => std_logic_vector'(x"00000000"),
  7116 => std_logic_vector'(x"00000000"),
  7117 => std_logic_vector'(x"00000000"),
  7118 => std_logic_vector'(x"00000000"),
  7119 => std_logic_vector'(x"00000000"),
  7120 => std_logic_vector'(x"00000000"),
  7121 => std_logic_vector'(x"00000000"),
  7122 => std_logic_vector'(x"00000000"),
  7123 => std_logic_vector'(x"00000000"),
  7124 => std_logic_vector'(x"00000000"),
  7125 => std_logic_vector'(x"00000000"),
  7126 => std_logic_vector'(x"00000000"),
  7127 => std_logic_vector'(x"00000000"),
  7128 => std_logic_vector'(x"00000000"),
  7129 => std_logic_vector'(x"00000000"),
  7130 => std_logic_vector'(x"00000000"),
  7131 => std_logic_vector'(x"00000000"),
  7132 => std_logic_vector'(x"00000000"),
  7133 => std_logic_vector'(x"00000000"),
  7134 => std_logic_vector'(x"00000000"),
  7135 => std_logic_vector'(x"00000000"),
  7136 => std_logic_vector'(x"00000000"),
  7137 => std_logic_vector'(x"00000000"),
  7138 => std_logic_vector'(x"00000000"),
  7139 => std_logic_vector'(x"00000000"),
  7140 => std_logic_vector'(x"00000000"),
  7141 => std_logic_vector'(x"00000000"),
  7142 => std_logic_vector'(x"00000000"),
  7143 => std_logic_vector'(x"00000000"),
  7144 => std_logic_vector'(x"00000000"),
  7145 => std_logic_vector'(x"00000000"),
  7146 => std_logic_vector'(x"00000000"),
  7147 => std_logic_vector'(x"00000000"),
  7148 => std_logic_vector'(x"00000000"),
  7149 => std_logic_vector'(x"00000000"),
  7150 => std_logic_vector'(x"00000000"),
  7151 => std_logic_vector'(x"00000000"),
  7152 => std_logic_vector'(x"00000000"),
  7153 => std_logic_vector'(x"00000000"),
  7154 => std_logic_vector'(x"00000000"),
  7155 => std_logic_vector'(x"00000000"),
  7156 => std_logic_vector'(x"00000000"),
  7157 => std_logic_vector'(x"00000000"),
  7158 => std_logic_vector'(x"00000000"),
  7159 => std_logic_vector'(x"00000000"),
  7160 => std_logic_vector'(x"00000000"),
  7161 => std_logic_vector'(x"00000000"),
  7162 => std_logic_vector'(x"00000000"),
  7163 => std_logic_vector'(x"00000000"),
  7164 => std_logic_vector'(x"00000000"),
  7165 => std_logic_vector'(x"00000000"),
  7166 => std_logic_vector'(x"00000000"),
  7167 => std_logic_vector'(x"00000000"),
  7168 => std_logic_vector'(x"00000000"),
  7169 => std_logic_vector'(x"00000000"),
  7170 => std_logic_vector'(x"00000000"),
  7171 => std_logic_vector'(x"00000000"),
  7172 => std_logic_vector'(x"00000000"),
  7173 => std_logic_vector'(x"00000000"),
  7174 => std_logic_vector'(x"00000000"),
  7175 => std_logic_vector'(x"00000000"),
  7176 => std_logic_vector'(x"00000000"),
  7177 => std_logic_vector'(x"00000000"),
  7178 => std_logic_vector'(x"00000000"),
  7179 => std_logic_vector'(x"00000000"),
  7180 => std_logic_vector'(x"00000000"),
  7181 => std_logic_vector'(x"00000000"),
  7182 => std_logic_vector'(x"00000000"),
  7183 => std_logic_vector'(x"00000000"),
  7184 => std_logic_vector'(x"00000000"),
  7185 => std_logic_vector'(x"00000000"),
  7186 => std_logic_vector'(x"00000000"),
  7187 => std_logic_vector'(x"00000000"),
  7188 => std_logic_vector'(x"00000000"),
  7189 => std_logic_vector'(x"00000000"),
  7190 => std_logic_vector'(x"00000000"),
  7191 => std_logic_vector'(x"00000000"),
  7192 => std_logic_vector'(x"00000000"),
  7193 => std_logic_vector'(x"00000000"),
  7194 => std_logic_vector'(x"00000000"),
  7195 => std_logic_vector'(x"00000000"),
  7196 => std_logic_vector'(x"00000000"),
  7197 => std_logic_vector'(x"00000000"),
  7198 => std_logic_vector'(x"00000000"),
  7199 => std_logic_vector'(x"00000000"),
  7200 => std_logic_vector'(x"00000000"),
  7201 => std_logic_vector'(x"00000000"),
  7202 => std_logic_vector'(x"00000000"),
  7203 => std_logic_vector'(x"00000000"),
  7204 => std_logic_vector'(x"00000000"),
  7205 => std_logic_vector'(x"00000000"),
  7206 => std_logic_vector'(x"00000000"),
  7207 => std_logic_vector'(x"00000000"),
  7208 => std_logic_vector'(x"00000000"),
  7209 => std_logic_vector'(x"00000000"),
  7210 => std_logic_vector'(x"00000000"),
  7211 => std_logic_vector'(x"00000000"),
  7212 => std_logic_vector'(x"00000000"),
  7213 => std_logic_vector'(x"00000000"),
  7214 => std_logic_vector'(x"00000000"),
  7215 => std_logic_vector'(x"00000000"),
  7216 => std_logic_vector'(x"00000000"),
  7217 => std_logic_vector'(x"00000000"),
  7218 => std_logic_vector'(x"00000000"),
  7219 => std_logic_vector'(x"00000000"),
  7220 => std_logic_vector'(x"00000000"),
  7221 => std_logic_vector'(x"00000000"),
  7222 => std_logic_vector'(x"00000000"),
  7223 => std_logic_vector'(x"00000000"),
  7224 => std_logic_vector'(x"00000000"),
  7225 => std_logic_vector'(x"00000000"),
  7226 => std_logic_vector'(x"00000000"),
  7227 => std_logic_vector'(x"00000000"),
  7228 => std_logic_vector'(x"00000000"),
  7229 => std_logic_vector'(x"00000000"),
  7230 => std_logic_vector'(x"00000000"),
  7231 => std_logic_vector'(x"00000000"),
  7232 => std_logic_vector'(x"00000000"),
  7233 => std_logic_vector'(x"00000000"),
  7234 => std_logic_vector'(x"00000000"),
  7235 => std_logic_vector'(x"00000000"),
  7236 => std_logic_vector'(x"00000000"),
  7237 => std_logic_vector'(x"00000000"),
  7238 => std_logic_vector'(x"00000000"),
  7239 => std_logic_vector'(x"00000000"),
  7240 => std_logic_vector'(x"00000000"),
  7241 => std_logic_vector'(x"00000000"),
  7242 => std_logic_vector'(x"00000000"),
  7243 => std_logic_vector'(x"00000000"),
  7244 => std_logic_vector'(x"00000000"),
  7245 => std_logic_vector'(x"00000000"),
  7246 => std_logic_vector'(x"00000000"),
  7247 => std_logic_vector'(x"00000000"),
  7248 => std_logic_vector'(x"00000000"),
  7249 => std_logic_vector'(x"00000000"),
  7250 => std_logic_vector'(x"00000000"),
  7251 => std_logic_vector'(x"00000000"),
  7252 => std_logic_vector'(x"00000000"),
  7253 => std_logic_vector'(x"00000000"),
  7254 => std_logic_vector'(x"00000000"),
  7255 => std_logic_vector'(x"00000000"),
  7256 => std_logic_vector'(x"00000000"),
  7257 => std_logic_vector'(x"00000000"),
  7258 => std_logic_vector'(x"00000000"),
  7259 => std_logic_vector'(x"00000000"),
  7260 => std_logic_vector'(x"00000000"),
  7261 => std_logic_vector'(x"00000000"),
  7262 => std_logic_vector'(x"00000000"),
  7263 => std_logic_vector'(x"00000000"),
  7264 => std_logic_vector'(x"00000000"),
  7265 => std_logic_vector'(x"00000000"),
  7266 => std_logic_vector'(x"00000000"),
  7267 => std_logic_vector'(x"00000000"),
  7268 => std_logic_vector'(x"00000000"),
  7269 => std_logic_vector'(x"00000000"),
  7270 => std_logic_vector'(x"00000000"),
  7271 => std_logic_vector'(x"00000000"),
  7272 => std_logic_vector'(x"00000000"),
  7273 => std_logic_vector'(x"00000000"),
  7274 => std_logic_vector'(x"00000000"),
  7275 => std_logic_vector'(x"00000000"),
  7276 => std_logic_vector'(x"00000000"),
  7277 => std_logic_vector'(x"00000000"),
  7278 => std_logic_vector'(x"00000000"),
  7279 => std_logic_vector'(x"00000000"),
  7280 => std_logic_vector'(x"00000000"),
  7281 => std_logic_vector'(x"00000000"),
  7282 => std_logic_vector'(x"00000000"),
  7283 => std_logic_vector'(x"00000000"),
  7284 => std_logic_vector'(x"00000000"),
  7285 => std_logic_vector'(x"00000000"),
  7286 => std_logic_vector'(x"00000000"),
  7287 => std_logic_vector'(x"00000000"),
  7288 => std_logic_vector'(x"00000000"),
  7289 => std_logic_vector'(x"00000000"),
  7290 => std_logic_vector'(x"00000000"),
  7291 => std_logic_vector'(x"00000000"),
  7292 => std_logic_vector'(x"00000000"),
  7293 => std_logic_vector'(x"00000000"),
  7294 => std_logic_vector'(x"00000000"),
  7295 => std_logic_vector'(x"00000000"),
  7296 => std_logic_vector'(x"00000000"),
  7297 => std_logic_vector'(x"00000000"),
  7298 => std_logic_vector'(x"00000000"),
  7299 => std_logic_vector'(x"00000000"),
  7300 => std_logic_vector'(x"00000000"),
  7301 => std_logic_vector'(x"00000000"),
  7302 => std_logic_vector'(x"00000000"),
  7303 => std_logic_vector'(x"00000000"),
  7304 => std_logic_vector'(x"00000000"),
  7305 => std_logic_vector'(x"00000000"),
  7306 => std_logic_vector'(x"00000000"),
  7307 => std_logic_vector'(x"00000000"),
  7308 => std_logic_vector'(x"00000000"),
  7309 => std_logic_vector'(x"00000000"),
  7310 => std_logic_vector'(x"00000000"),
  7311 => std_logic_vector'(x"00000000"),
  7312 => std_logic_vector'(x"00000000"),
  7313 => std_logic_vector'(x"00000000"),
  7314 => std_logic_vector'(x"00000000"),
  7315 => std_logic_vector'(x"00000000"),
  7316 => std_logic_vector'(x"00000000"),
  7317 => std_logic_vector'(x"00000000"),
  7318 => std_logic_vector'(x"00000000"),
  7319 => std_logic_vector'(x"00000000"),
  7320 => std_logic_vector'(x"00000000"),
  7321 => std_logic_vector'(x"00000000"),
  7322 => std_logic_vector'(x"00000000"),
  7323 => std_logic_vector'(x"00000000"),
  7324 => std_logic_vector'(x"00000000"),
  7325 => std_logic_vector'(x"00000000"),
  7326 => std_logic_vector'(x"00000000"),
  7327 => std_logic_vector'(x"00000000"),
  7328 => std_logic_vector'(x"00000000"),
  7329 => std_logic_vector'(x"00000000"),
  7330 => std_logic_vector'(x"00000000"),
  7331 => std_logic_vector'(x"00000000"),
  7332 => std_logic_vector'(x"00000000"),
  7333 => std_logic_vector'(x"00000000"),
  7334 => std_logic_vector'(x"00000000"),
  7335 => std_logic_vector'(x"00000000"),
  7336 => std_logic_vector'(x"00000000"),
  7337 => std_logic_vector'(x"00000000"),
  7338 => std_logic_vector'(x"00000000"),
  7339 => std_logic_vector'(x"00000000"),
  7340 => std_logic_vector'(x"00000000"),
  7341 => std_logic_vector'(x"00000000"),
  7342 => std_logic_vector'(x"00000000"),
  7343 => std_logic_vector'(x"00000000"),
  7344 => std_logic_vector'(x"00000000"),
  7345 => std_logic_vector'(x"00000000"),
  7346 => std_logic_vector'(x"00000000"),
  7347 => std_logic_vector'(x"00000000"),
  7348 => std_logic_vector'(x"00000000"),
  7349 => std_logic_vector'(x"00000000"),
  7350 => std_logic_vector'(x"00000000"),
  7351 => std_logic_vector'(x"00000000"),
  7352 => std_logic_vector'(x"00000000"),
  7353 => std_logic_vector'(x"00000000"),
  7354 => std_logic_vector'(x"00000000"),
  7355 => std_logic_vector'(x"00000000"),
  7356 => std_logic_vector'(x"00000000"),
  7357 => std_logic_vector'(x"00000000"),
  7358 => std_logic_vector'(x"00000000"),
  7359 => std_logic_vector'(x"00000000"),
  7360 => std_logic_vector'(x"00000000"),
  7361 => std_logic_vector'(x"00000000"),
  7362 => std_logic_vector'(x"00000000"),
  7363 => std_logic_vector'(x"00000000"),
  7364 => std_logic_vector'(x"00000000"),
  7365 => std_logic_vector'(x"00000000"),
  7366 => std_logic_vector'(x"00000000"),
  7367 => std_logic_vector'(x"00000000"),
  7368 => std_logic_vector'(x"00000000"),
  7369 => std_logic_vector'(x"00000000"),
  7370 => std_logic_vector'(x"00000000"),
  7371 => std_logic_vector'(x"00000000"),
  7372 => std_logic_vector'(x"00000000"),
  7373 => std_logic_vector'(x"00000000"),
  7374 => std_logic_vector'(x"00000000"),
  7375 => std_logic_vector'(x"00000000"),
  7376 => std_logic_vector'(x"00000000"),
  7377 => std_logic_vector'(x"00000000"),
  7378 => std_logic_vector'(x"00000000"),
  7379 => std_logic_vector'(x"00000000"),
  7380 => std_logic_vector'(x"00000000"),
  7381 => std_logic_vector'(x"00000000"),
  7382 => std_logic_vector'(x"00000000"),
  7383 => std_logic_vector'(x"00000000"),
  7384 => std_logic_vector'(x"00000000"),
  7385 => std_logic_vector'(x"00000000"),
  7386 => std_logic_vector'(x"00000000"),
  7387 => std_logic_vector'(x"00000000"),
  7388 => std_logic_vector'(x"00000000"),
  7389 => std_logic_vector'(x"00000000"),
  7390 => std_logic_vector'(x"00000000"),
  7391 => std_logic_vector'(x"00000000"),
  7392 => std_logic_vector'(x"00000000"),
  7393 => std_logic_vector'(x"00000000"),
  7394 => std_logic_vector'(x"00000000"),
  7395 => std_logic_vector'(x"00000000"),
  7396 => std_logic_vector'(x"00000000"),
  7397 => std_logic_vector'(x"00000000"),
  7398 => std_logic_vector'(x"00000000"),
  7399 => std_logic_vector'(x"00000000"),
  7400 => std_logic_vector'(x"00000000"),
  7401 => std_logic_vector'(x"00000000"),
  7402 => std_logic_vector'(x"00000000"),
  7403 => std_logic_vector'(x"00000000"),
  7404 => std_logic_vector'(x"00000000"),
  7405 => std_logic_vector'(x"00000000"),
  7406 => std_logic_vector'(x"00000000"),
  7407 => std_logic_vector'(x"00000000"),
  7408 => std_logic_vector'(x"00000000"),
  7409 => std_logic_vector'(x"00000000"),
  7410 => std_logic_vector'(x"00000000"),
  7411 => std_logic_vector'(x"00000000"),
  7412 => std_logic_vector'(x"00000000"),
  7413 => std_logic_vector'(x"00000000"),
  7414 => std_logic_vector'(x"00000000"),
  7415 => std_logic_vector'(x"00000000"),
  7416 => std_logic_vector'(x"00000000"),
  7417 => std_logic_vector'(x"00000000"),
  7418 => std_logic_vector'(x"00000000"),
  7419 => std_logic_vector'(x"00000000"),
  7420 => std_logic_vector'(x"00000000"),
  7421 => std_logic_vector'(x"00000000"),
  7422 => std_logic_vector'(x"00000000"),
  7423 => std_logic_vector'(x"00000000"),
  7424 => std_logic_vector'(x"00000000"),
  7425 => std_logic_vector'(x"00000000"),
  7426 => std_logic_vector'(x"00000000"),
  7427 => std_logic_vector'(x"00000000"),
  7428 => std_logic_vector'(x"00000000"),
  7429 => std_logic_vector'(x"00000000"),
  7430 => std_logic_vector'(x"00000000"),
  7431 => std_logic_vector'(x"00000000"),
  7432 => std_logic_vector'(x"00000000"),
  7433 => std_logic_vector'(x"00000000"),
  7434 => std_logic_vector'(x"00000000"),
  7435 => std_logic_vector'(x"00000000"),
  7436 => std_logic_vector'(x"00000000"),
  7437 => std_logic_vector'(x"00000000"),
  7438 => std_logic_vector'(x"00000000"),
  7439 => std_logic_vector'(x"00000000"),
  7440 => std_logic_vector'(x"00000000"),
  7441 => std_logic_vector'(x"00000000"),
  7442 => std_logic_vector'(x"00000000"),
  7443 => std_logic_vector'(x"00000000"),
  7444 => std_logic_vector'(x"00000000"),
  7445 => std_logic_vector'(x"00000000"),
  7446 => std_logic_vector'(x"00000000"),
  7447 => std_logic_vector'(x"00000000"),
  7448 => std_logic_vector'(x"00000000"),
  7449 => std_logic_vector'(x"00000000"),
  7450 => std_logic_vector'(x"00000000"),
  7451 => std_logic_vector'(x"00000000"),
  7452 => std_logic_vector'(x"00000000"),
  7453 => std_logic_vector'(x"00000000"),
  7454 => std_logic_vector'(x"00000000"),
  7455 => std_logic_vector'(x"00000000"),
  7456 => std_logic_vector'(x"00000000"),
  7457 => std_logic_vector'(x"00000000"),
  7458 => std_logic_vector'(x"00000000"),
  7459 => std_logic_vector'(x"00000000"),
  7460 => std_logic_vector'(x"00000000"),
  7461 => std_logic_vector'(x"00000000"),
  7462 => std_logic_vector'(x"00000000"),
  7463 => std_logic_vector'(x"00000000"),
  7464 => std_logic_vector'(x"00000000"),
  7465 => std_logic_vector'(x"00000000"),
  7466 => std_logic_vector'(x"00000000"),
  7467 => std_logic_vector'(x"00000000"),
  7468 => std_logic_vector'(x"00000000"),
  7469 => std_logic_vector'(x"00000000"),
  7470 => std_logic_vector'(x"00000000"),
  7471 => std_logic_vector'(x"00000000"),
  7472 => std_logic_vector'(x"00000000"),
  7473 => std_logic_vector'(x"00000000"),
  7474 => std_logic_vector'(x"00000000"),
  7475 => std_logic_vector'(x"00000000"),
  7476 => std_logic_vector'(x"00000000"),
  7477 => std_logic_vector'(x"00000000"),
  7478 => std_logic_vector'(x"00000000"),
  7479 => std_logic_vector'(x"00000000"),
  7480 => std_logic_vector'(x"00000000"),
  7481 => std_logic_vector'(x"00000000"),
  7482 => std_logic_vector'(x"00000000"),
  7483 => std_logic_vector'(x"00000000"),
  7484 => std_logic_vector'(x"00000000"),
  7485 => std_logic_vector'(x"00000000"),
  7486 => std_logic_vector'(x"00000000"),
  7487 => std_logic_vector'(x"00000000"),
  7488 => std_logic_vector'(x"00000000"),
  7489 => std_logic_vector'(x"00000000"),
  7490 => std_logic_vector'(x"00000000"),
  7491 => std_logic_vector'(x"00000000"),
  7492 => std_logic_vector'(x"00000000"),
  7493 => std_logic_vector'(x"00000000"),
  7494 => std_logic_vector'(x"00000000"),
  7495 => std_logic_vector'(x"00000000"),
  7496 => std_logic_vector'(x"00000000"),
  7497 => std_logic_vector'(x"00000000"),
  7498 => std_logic_vector'(x"00000000"),
  7499 => std_logic_vector'(x"00000000"),
  7500 => std_logic_vector'(x"00000000"),
  7501 => std_logic_vector'(x"00000000"),
  7502 => std_logic_vector'(x"00000000"),
  7503 => std_logic_vector'(x"00000000"),
  7504 => std_logic_vector'(x"00000000"),
  7505 => std_logic_vector'(x"00000000"),
  7506 => std_logic_vector'(x"00000000"),
  7507 => std_logic_vector'(x"00000000"),
  7508 => std_logic_vector'(x"00000000"),
  7509 => std_logic_vector'(x"00000000"),
  7510 => std_logic_vector'(x"00000000"),
  7511 => std_logic_vector'(x"00000000"),
  7512 => std_logic_vector'(x"00000000"),
  7513 => std_logic_vector'(x"00000000"),
  7514 => std_logic_vector'(x"00000000"),
  7515 => std_logic_vector'(x"00000000"),
  7516 => std_logic_vector'(x"00000000"),
  7517 => std_logic_vector'(x"00000000"),
  7518 => std_logic_vector'(x"00000000"),
  7519 => std_logic_vector'(x"00000000"),
  7520 => std_logic_vector'(x"00000000"),
  7521 => std_logic_vector'(x"00000000"),
  7522 => std_logic_vector'(x"00000000"),
  7523 => std_logic_vector'(x"00000000"),
  7524 => std_logic_vector'(x"00000000"),
  7525 => std_logic_vector'(x"00000000"),
  7526 => std_logic_vector'(x"00000000"),
  7527 => std_logic_vector'(x"00000000"),
  7528 => std_logic_vector'(x"00000000"),
  7529 => std_logic_vector'(x"00000000"),
  7530 => std_logic_vector'(x"00000000"),
  7531 => std_logic_vector'(x"00000000"),
  7532 => std_logic_vector'(x"00000000"),
  7533 => std_logic_vector'(x"00000000"),
  7534 => std_logic_vector'(x"00000000"),
  7535 => std_logic_vector'(x"00000000"),
  7536 => std_logic_vector'(x"00000000"),
  7537 => std_logic_vector'(x"00000000"),
  7538 => std_logic_vector'(x"00000000"),
  7539 => std_logic_vector'(x"00000000"),
  7540 => std_logic_vector'(x"00000000"),
  7541 => std_logic_vector'(x"00000000"),
  7542 => std_logic_vector'(x"00000000"),
  7543 => std_logic_vector'(x"00000000"),
  7544 => std_logic_vector'(x"00000000"),
  7545 => std_logic_vector'(x"00000000"),
  7546 => std_logic_vector'(x"00000000"),
  7547 => std_logic_vector'(x"00000000"),
  7548 => std_logic_vector'(x"00000000"),
  7549 => std_logic_vector'(x"00000000"),
  7550 => std_logic_vector'(x"00000000"),
  7551 => std_logic_vector'(x"00000000"),
  7552 => std_logic_vector'(x"00000000"),
  7553 => std_logic_vector'(x"00000000"),
  7554 => std_logic_vector'(x"00000000"),
  7555 => std_logic_vector'(x"00000000"),
  7556 => std_logic_vector'(x"00000000"),
  7557 => std_logic_vector'(x"00000000"),
  7558 => std_logic_vector'(x"00000000"),
  7559 => std_logic_vector'(x"00000000"),
  7560 => std_logic_vector'(x"00000000"),
  7561 => std_logic_vector'(x"00000000"),
  7562 => std_logic_vector'(x"00000000"),
  7563 => std_logic_vector'(x"00000000"),
  7564 => std_logic_vector'(x"00000000"),
  7565 => std_logic_vector'(x"00000000"),
  7566 => std_logic_vector'(x"00000000"),
  7567 => std_logic_vector'(x"00000000"),
  7568 => std_logic_vector'(x"00000000"),
  7569 => std_logic_vector'(x"00000000"),
  7570 => std_logic_vector'(x"00000000"),
  7571 => std_logic_vector'(x"00000000"),
  7572 => std_logic_vector'(x"00000000"),
  7573 => std_logic_vector'(x"00000000"),
  7574 => std_logic_vector'(x"00000000"),
  7575 => std_logic_vector'(x"00000000"),
  7576 => std_logic_vector'(x"00000000"),
  7577 => std_logic_vector'(x"00000000"),
  7578 => std_logic_vector'(x"00000000"),
  7579 => std_logic_vector'(x"00000000"),
  7580 => std_logic_vector'(x"00000000"),
  7581 => std_logic_vector'(x"00000000"),
  7582 => std_logic_vector'(x"00000000"),
  7583 => std_logic_vector'(x"00000000"),
  7584 => std_logic_vector'(x"00000000"),
  7585 => std_logic_vector'(x"00000000"),
  7586 => std_logic_vector'(x"00000000"),
  7587 => std_logic_vector'(x"00000000"),
  7588 => std_logic_vector'(x"00000000"),
  7589 => std_logic_vector'(x"00000000"),
  7590 => std_logic_vector'(x"00000000"),
  7591 => std_logic_vector'(x"00000000"),
  7592 => std_logic_vector'(x"00000000"),
  7593 => std_logic_vector'(x"00000000"),
  7594 => std_logic_vector'(x"00000000"),
  7595 => std_logic_vector'(x"00000000"),
  7596 => std_logic_vector'(x"00000000"),
  7597 => std_logic_vector'(x"00000000"),
  7598 => std_logic_vector'(x"00000000"),
  7599 => std_logic_vector'(x"00000000"),
  7600 => std_logic_vector'(x"00000000"),
  7601 => std_logic_vector'(x"00000000"),
  7602 => std_logic_vector'(x"00000000"),
  7603 => std_logic_vector'(x"00000000"),
  7604 => std_logic_vector'(x"00000000"),
  7605 => std_logic_vector'(x"00000000"),
  7606 => std_logic_vector'(x"00000000"),
  7607 => std_logic_vector'(x"00000000"),
  7608 => std_logic_vector'(x"00000000"),
  7609 => std_logic_vector'(x"00000000"),
  7610 => std_logic_vector'(x"00000000"),
  7611 => std_logic_vector'(x"00000000"),
  7612 => std_logic_vector'(x"00000000"),
  7613 => std_logic_vector'(x"00000000"),
  7614 => std_logic_vector'(x"00000000"),
  7615 => std_logic_vector'(x"00000000"),
  7616 => std_logic_vector'(x"00000000"),
  7617 => std_logic_vector'(x"00000000"),
  7618 => std_logic_vector'(x"00000000"),
  7619 => std_logic_vector'(x"00000000"),
  7620 => std_logic_vector'(x"00000000"),
  7621 => std_logic_vector'(x"00000000"),
  7622 => std_logic_vector'(x"00000000"),
  7623 => std_logic_vector'(x"00000000"),
  7624 => std_logic_vector'(x"00000000"),
  7625 => std_logic_vector'(x"00000000"),
  7626 => std_logic_vector'(x"00000000"),
  7627 => std_logic_vector'(x"00000000"),
  7628 => std_logic_vector'(x"00000000"),
  7629 => std_logic_vector'(x"00000000"),
  7630 => std_logic_vector'(x"00000000"),
  7631 => std_logic_vector'(x"00000000"),
  7632 => std_logic_vector'(x"00000000"),
  7633 => std_logic_vector'(x"00000000"),
  7634 => std_logic_vector'(x"00000000"),
  7635 => std_logic_vector'(x"00000000"),
  7636 => std_logic_vector'(x"00000000"),
  7637 => std_logic_vector'(x"00000000"),
  7638 => std_logic_vector'(x"00000000"),
  7639 => std_logic_vector'(x"00000000"),
  7640 => std_logic_vector'(x"00000000"),
  7641 => std_logic_vector'(x"00000000"),
  7642 => std_logic_vector'(x"00000000"),
  7643 => std_logic_vector'(x"00000000"),
  7644 => std_logic_vector'(x"00000000"),
  7645 => std_logic_vector'(x"00000000"),
  7646 => std_logic_vector'(x"00000000"),
  7647 => std_logic_vector'(x"00000000"),
  7648 => std_logic_vector'(x"00000000"),
  7649 => std_logic_vector'(x"00000000"),
  7650 => std_logic_vector'(x"00000000"),
  7651 => std_logic_vector'(x"00000000"),
  7652 => std_logic_vector'(x"00000000"),
  7653 => std_logic_vector'(x"00000000"),
  7654 => std_logic_vector'(x"00000000"),
  7655 => std_logic_vector'(x"00000000"),
  7656 => std_logic_vector'(x"00000000"),
  7657 => std_logic_vector'(x"00000000"),
  7658 => std_logic_vector'(x"00000000"),
  7659 => std_logic_vector'(x"00000000"),
  7660 => std_logic_vector'(x"00000000"),
  7661 => std_logic_vector'(x"00000000"),
  7662 => std_logic_vector'(x"00000000"),
  7663 => std_logic_vector'(x"00000000"),
  7664 => std_logic_vector'(x"00000000"),
  7665 => std_logic_vector'(x"00000000"),
  7666 => std_logic_vector'(x"00000000"),
  7667 => std_logic_vector'(x"00000000"),
  7668 => std_logic_vector'(x"00000000"),
  7669 => std_logic_vector'(x"00000000"),
  7670 => std_logic_vector'(x"00000000"),
  7671 => std_logic_vector'(x"00000000"),
  7672 => std_logic_vector'(x"00000000"),
  7673 => std_logic_vector'(x"00000000"),
  7674 => std_logic_vector'(x"00000000"),
  7675 => std_logic_vector'(x"00000000"),
  7676 => std_logic_vector'(x"00000000"),
  7677 => std_logic_vector'(x"00000000"),
  7678 => std_logic_vector'(x"00000000"),
  7679 => std_logic_vector'(x"00000000"),
  7680 => std_logic_vector'(x"00000000"),
  7681 => std_logic_vector'(x"00000000"),
  7682 => std_logic_vector'(x"00000000"),
  7683 => std_logic_vector'(x"00000000"),
  7684 => std_logic_vector'(x"00000000"),
  7685 => std_logic_vector'(x"00000000"),
  7686 => std_logic_vector'(x"00000000"),
  7687 => std_logic_vector'(x"00000000"),
  7688 => std_logic_vector'(x"00000000"),
  7689 => std_logic_vector'(x"00000000"),
  7690 => std_logic_vector'(x"00000000"),
  7691 => std_logic_vector'(x"00000000"),
  7692 => std_logic_vector'(x"00000000"),
  7693 => std_logic_vector'(x"00000000"),
  7694 => std_logic_vector'(x"00000000"),
  7695 => std_logic_vector'(x"00000000"),
  7696 => std_logic_vector'(x"00000000"),
  7697 => std_logic_vector'(x"00000000"),
  7698 => std_logic_vector'(x"00000000"),
  7699 => std_logic_vector'(x"00000000"),
  7700 => std_logic_vector'(x"00000000"),
  7701 => std_logic_vector'(x"00000000"),
  7702 => std_logic_vector'(x"00000000"),
  7703 => std_logic_vector'(x"00000000"),
  7704 => std_logic_vector'(x"00000000"),
  7705 => std_logic_vector'(x"00000000"),
  7706 => std_logic_vector'(x"00000000"),
  7707 => std_logic_vector'(x"00000000"),
  7708 => std_logic_vector'(x"00000000"),
  7709 => std_logic_vector'(x"00000000"),
  7710 => std_logic_vector'(x"00000000"),
  7711 => std_logic_vector'(x"00000000"),
  7712 => std_logic_vector'(x"00000000"),
  7713 => std_logic_vector'(x"00000000"),
  7714 => std_logic_vector'(x"00000000"),
  7715 => std_logic_vector'(x"00000000"),
  7716 => std_logic_vector'(x"00000000"),
  7717 => std_logic_vector'(x"00000000"),
  7718 => std_logic_vector'(x"00000000"),
  7719 => std_logic_vector'(x"00000000"),
  7720 => std_logic_vector'(x"00000000"),
  7721 => std_logic_vector'(x"00000000"),
  7722 => std_logic_vector'(x"00000000"),
  7723 => std_logic_vector'(x"00000000"),
  7724 => std_logic_vector'(x"00000000"),
  7725 => std_logic_vector'(x"00000000"),
  7726 => std_logic_vector'(x"00000000"),
  7727 => std_logic_vector'(x"00000000"),
  7728 => std_logic_vector'(x"00000000"),
  7729 => std_logic_vector'(x"00000000"),
  7730 => std_logic_vector'(x"00000000"),
  7731 => std_logic_vector'(x"00000000"),
  7732 => std_logic_vector'(x"00000000"),
  7733 => std_logic_vector'(x"00000000"),
  7734 => std_logic_vector'(x"00000000"),
  7735 => std_logic_vector'(x"00000000"),
  7736 => std_logic_vector'(x"00000000"),
  7737 => std_logic_vector'(x"00000000"),
  7738 => std_logic_vector'(x"00000000"),
  7739 => std_logic_vector'(x"00000000"),
  7740 => std_logic_vector'(x"00000000"),
  7741 => std_logic_vector'(x"00000000"),
  7742 => std_logic_vector'(x"00000000"),
  7743 => std_logic_vector'(x"00000000"),
  7744 => std_logic_vector'(x"00000000"),
  7745 => std_logic_vector'(x"00000000"),
  7746 => std_logic_vector'(x"00000000"),
  7747 => std_logic_vector'(x"00000000"),
  7748 => std_logic_vector'(x"00000000"),
  7749 => std_logic_vector'(x"00000000"),
  7750 => std_logic_vector'(x"00000000"),
  7751 => std_logic_vector'(x"00000000"),
  7752 => std_logic_vector'(x"00000000"),
  7753 => std_logic_vector'(x"00000000"),
  7754 => std_logic_vector'(x"00000000"),
  7755 => std_logic_vector'(x"00000000"),
  7756 => std_logic_vector'(x"00000000"),
  7757 => std_logic_vector'(x"00000000"),
  7758 => std_logic_vector'(x"00000000"),
  7759 => std_logic_vector'(x"00000000"),
  7760 => std_logic_vector'(x"00000000"),
  7761 => std_logic_vector'(x"00000000"),
  7762 => std_logic_vector'(x"00000000"),
  7763 => std_logic_vector'(x"00000000"),
  7764 => std_logic_vector'(x"00000000"),
  7765 => std_logic_vector'(x"00000000"),
  7766 => std_logic_vector'(x"00000000"),
  7767 => std_logic_vector'(x"00000000"),
  7768 => std_logic_vector'(x"00000000"),
  7769 => std_logic_vector'(x"00000000"),
  7770 => std_logic_vector'(x"00000000"),
  7771 => std_logic_vector'(x"00000000"),
  7772 => std_logic_vector'(x"00000000"),
  7773 => std_logic_vector'(x"00000000"),
  7774 => std_logic_vector'(x"00000000"),
  7775 => std_logic_vector'(x"00000000"),
  7776 => std_logic_vector'(x"00000000"),
  7777 => std_logic_vector'(x"00000000"),
  7778 => std_logic_vector'(x"00000000"),
  7779 => std_logic_vector'(x"00000000"),
  7780 => std_logic_vector'(x"00000000"),
  7781 => std_logic_vector'(x"00000000"),
  7782 => std_logic_vector'(x"00000000"),
  7783 => std_logic_vector'(x"00000000"),
  7784 => std_logic_vector'(x"00000000"),
  7785 => std_logic_vector'(x"00000000"),
  7786 => std_logic_vector'(x"00000000"),
  7787 => std_logic_vector'(x"00000000"),
  7788 => std_logic_vector'(x"00000000"),
  7789 => std_logic_vector'(x"00000000"),
  7790 => std_logic_vector'(x"00000000"),
  7791 => std_logic_vector'(x"00000000"),
  7792 => std_logic_vector'(x"00000000"),
  7793 => std_logic_vector'(x"00000000"),
  7794 => std_logic_vector'(x"00000000"),
  7795 => std_logic_vector'(x"00000000"),
  7796 => std_logic_vector'(x"00000000"),
  7797 => std_logic_vector'(x"00000000"),
  7798 => std_logic_vector'(x"00000000"),
  7799 => std_logic_vector'(x"00000000"),
  7800 => std_logic_vector'(x"00000000"),
  7801 => std_logic_vector'(x"00000000"),
  7802 => std_logic_vector'(x"00000000"),
  7803 => std_logic_vector'(x"00000000"),
  7804 => std_logic_vector'(x"00000000"),
  7805 => std_logic_vector'(x"00000000"),
  7806 => std_logic_vector'(x"00000000"),
  7807 => std_logic_vector'(x"00000000"),
  7808 => std_logic_vector'(x"00000000"),
  7809 => std_logic_vector'(x"00000000"),
  7810 => std_logic_vector'(x"00000000"),
  7811 => std_logic_vector'(x"00000000"),
  7812 => std_logic_vector'(x"00000000"),
  7813 => std_logic_vector'(x"00000000"),
  7814 => std_logic_vector'(x"00000000"),
  7815 => std_logic_vector'(x"00000000"),
  7816 => std_logic_vector'(x"00000000"),
  7817 => std_logic_vector'(x"00000000"),
  7818 => std_logic_vector'(x"00000000"),
  7819 => std_logic_vector'(x"00000000"),
  7820 => std_logic_vector'(x"00000000"),
  7821 => std_logic_vector'(x"00000000"),
  7822 => std_logic_vector'(x"00000000"),
  7823 => std_logic_vector'(x"00000000"),
  7824 => std_logic_vector'(x"00000000"),
  7825 => std_logic_vector'(x"00000000"),
  7826 => std_logic_vector'(x"00000000"),
  7827 => std_logic_vector'(x"00000000"),
  7828 => std_logic_vector'(x"00000000"),
  7829 => std_logic_vector'(x"00000000"),
  7830 => std_logic_vector'(x"00000000"),
  7831 => std_logic_vector'(x"00000000"),
  7832 => std_logic_vector'(x"00000000"),
  7833 => std_logic_vector'(x"00000000"),
  7834 => std_logic_vector'(x"00000000"),
  7835 => std_logic_vector'(x"00000000"),
  7836 => std_logic_vector'(x"00000000"),
  7837 => std_logic_vector'(x"00000000"),
  7838 => std_logic_vector'(x"00000000"),
  7839 => std_logic_vector'(x"00000000"),
  7840 => std_logic_vector'(x"00000000"),
  7841 => std_logic_vector'(x"00000000"),
  7842 => std_logic_vector'(x"00000000"),
  7843 => std_logic_vector'(x"00000000"),
  7844 => std_logic_vector'(x"00000000"),
  7845 => std_logic_vector'(x"00000000"),
  7846 => std_logic_vector'(x"00000000"),
  7847 => std_logic_vector'(x"00000000"),
  7848 => std_logic_vector'(x"00000000"),
  7849 => std_logic_vector'(x"00000000"),
  7850 => std_logic_vector'(x"00000000"),
  7851 => std_logic_vector'(x"00000000"),
  7852 => std_logic_vector'(x"00000000"),
  7853 => std_logic_vector'(x"00000000"),
  7854 => std_logic_vector'(x"00000000"),
  7855 => std_logic_vector'(x"00000000"),
  7856 => std_logic_vector'(x"00000000"),
  7857 => std_logic_vector'(x"00000000"),
  7858 => std_logic_vector'(x"00000000"),
  7859 => std_logic_vector'(x"00000000"),
  7860 => std_logic_vector'(x"00000000"),
  7861 => std_logic_vector'(x"00000000"),
  7862 => std_logic_vector'(x"00000000"),
  7863 => std_logic_vector'(x"00000000"),
  7864 => std_logic_vector'(x"00000000"),
  7865 => std_logic_vector'(x"00000000"),
  7866 => std_logic_vector'(x"00000000"),
  7867 => std_logic_vector'(x"00000000"),
  7868 => std_logic_vector'(x"00000000"),
  7869 => std_logic_vector'(x"00000000"),
  7870 => std_logic_vector'(x"00000000"),
  7871 => std_logic_vector'(x"00000000"),
  7872 => std_logic_vector'(x"00000000"),
  7873 => std_logic_vector'(x"00000000"),
  7874 => std_logic_vector'(x"00000000"),
  7875 => std_logic_vector'(x"00000000"),
  7876 => std_logic_vector'(x"00000000"),
  7877 => std_logic_vector'(x"00000000"),
  7878 => std_logic_vector'(x"00000000"),
  7879 => std_logic_vector'(x"00000000"),
  7880 => std_logic_vector'(x"00000000"),
  7881 => std_logic_vector'(x"00000000"),
  7882 => std_logic_vector'(x"00000000"),
  7883 => std_logic_vector'(x"00000000"),
  7884 => std_logic_vector'(x"00000000"),
  7885 => std_logic_vector'(x"00000000"),
  7886 => std_logic_vector'(x"00000000"),
  7887 => std_logic_vector'(x"00000000"),
  7888 => std_logic_vector'(x"00000000"),
  7889 => std_logic_vector'(x"00000000"),
  7890 => std_logic_vector'(x"00000000"),
  7891 => std_logic_vector'(x"00000000"),
  7892 => std_logic_vector'(x"00000000"),
  7893 => std_logic_vector'(x"00000000"),
  7894 => std_logic_vector'(x"00000000"),
  7895 => std_logic_vector'(x"00000000"),
  7896 => std_logic_vector'(x"00000000"),
  7897 => std_logic_vector'(x"00000000"),
  7898 => std_logic_vector'(x"00000000"),
  7899 => std_logic_vector'(x"00000000"),
  7900 => std_logic_vector'(x"00000000"),
  7901 => std_logic_vector'(x"00000000"),
  7902 => std_logic_vector'(x"00000000"),
  7903 => std_logic_vector'(x"00000000"),
  7904 => std_logic_vector'(x"00000000"),
  7905 => std_logic_vector'(x"00000000"),
  7906 => std_logic_vector'(x"00000000"),
  7907 => std_logic_vector'(x"00000000"),
  7908 => std_logic_vector'(x"00000000"),
  7909 => std_logic_vector'(x"00000000"),
  7910 => std_logic_vector'(x"00000000"),
  7911 => std_logic_vector'(x"00000000"),
  7912 => std_logic_vector'(x"00000000"),
  7913 => std_logic_vector'(x"00000000"),
  7914 => std_logic_vector'(x"00000000"),
  7915 => std_logic_vector'(x"00000000"),
  7916 => std_logic_vector'(x"00000000"),
  7917 => std_logic_vector'(x"00000000"),
  7918 => std_logic_vector'(x"00000000"),
  7919 => std_logic_vector'(x"00000000"),
  7920 => std_logic_vector'(x"00000000"),
  7921 => std_logic_vector'(x"00000000"),
  7922 => std_logic_vector'(x"00000000"),
  7923 => std_logic_vector'(x"00000000"),
  7924 => std_logic_vector'(x"00000000"),
  7925 => std_logic_vector'(x"00000000"),
  7926 => std_logic_vector'(x"00000000"),
  7927 => std_logic_vector'(x"00000000"),
  7928 => std_logic_vector'(x"00000000"),
  7929 => std_logic_vector'(x"00000000"),
  7930 => std_logic_vector'(x"00000000"),
  7931 => std_logic_vector'(x"00000000"),
  7932 => std_logic_vector'(x"00000000"),
  7933 => std_logic_vector'(x"00000000"),
  7934 => std_logic_vector'(x"00000000"),
  7935 => std_logic_vector'(x"00000000"),
  7936 => std_logic_vector'(x"00000000"),
  7937 => std_logic_vector'(x"00000000"),
  7938 => std_logic_vector'(x"00000000"),
  7939 => std_logic_vector'(x"00000000"),
  7940 => std_logic_vector'(x"00000000"),
  7941 => std_logic_vector'(x"00000000"),
  7942 => std_logic_vector'(x"00000000"),
  7943 => std_logic_vector'(x"00000000"),
  7944 => std_logic_vector'(x"00000000"),
  7945 => std_logic_vector'(x"00000000"),
  7946 => std_logic_vector'(x"00000000"),
  7947 => std_logic_vector'(x"00000000"),
  7948 => std_logic_vector'(x"00000000"),
  7949 => std_logic_vector'(x"00000000"),
  7950 => std_logic_vector'(x"00000000"),
  7951 => std_logic_vector'(x"00000000"),
  7952 => std_logic_vector'(x"00000000"),
  7953 => std_logic_vector'(x"00000000"),
  7954 => std_logic_vector'(x"00000000"),
  7955 => std_logic_vector'(x"00000000"),
  7956 => std_logic_vector'(x"00000000"),
  7957 => std_logic_vector'(x"00000000"),
  7958 => std_logic_vector'(x"00000000"),
  7959 => std_logic_vector'(x"00000000"),
  7960 => std_logic_vector'(x"00000000"),
  7961 => std_logic_vector'(x"00000000"),
  7962 => std_logic_vector'(x"00000000"),
  7963 => std_logic_vector'(x"00000000"),
  7964 => std_logic_vector'(x"00000000"),
  7965 => std_logic_vector'(x"00000000"),
  7966 => std_logic_vector'(x"00000000"),
  7967 => std_logic_vector'(x"00000000"),
  7968 => std_logic_vector'(x"00000000"),
  7969 => std_logic_vector'(x"00000000"),
  7970 => std_logic_vector'(x"00000000"),
  7971 => std_logic_vector'(x"00000000"),
  7972 => std_logic_vector'(x"00000000"),
  7973 => std_logic_vector'(x"00000000"),
  7974 => std_logic_vector'(x"00000000"),
  7975 => std_logic_vector'(x"00000000"),
  7976 => std_logic_vector'(x"00000000"),
  7977 => std_logic_vector'(x"00000000"),
  7978 => std_logic_vector'(x"00000000"),
  7979 => std_logic_vector'(x"00000000"),
  7980 => std_logic_vector'(x"00000000"),
  7981 => std_logic_vector'(x"00000000"),
  7982 => std_logic_vector'(x"00000000"),
  7983 => std_logic_vector'(x"00000000"),
  7984 => std_logic_vector'(x"00000000"),
  7985 => std_logic_vector'(x"00000000"),
  7986 => std_logic_vector'(x"00000000"),
  7987 => std_logic_vector'(x"00000000"),
  7988 => std_logic_vector'(x"00000000"),
  7989 => std_logic_vector'(x"00000000"),
  7990 => std_logic_vector'(x"00000000"),
  7991 => std_logic_vector'(x"00000000"),
  7992 => std_logic_vector'(x"00000000"),
  7993 => std_logic_vector'(x"00000000"),
  7994 => std_logic_vector'(x"00000000"),
  7995 => std_logic_vector'(x"00000000"),
  7996 => std_logic_vector'(x"00000000"),
  7997 => std_logic_vector'(x"00000000"),
  7998 => std_logic_vector'(x"00000000"),
  7999 => std_logic_vector'(x"00000000"),
  8000 => std_logic_vector'(x"00000000"),
  8001 => std_logic_vector'(x"00000000"),
  8002 => std_logic_vector'(x"00000000"),
  8003 => std_logic_vector'(x"00000000"),
  8004 => std_logic_vector'(x"00000000"),
  8005 => std_logic_vector'(x"00000000"),
  8006 => std_logic_vector'(x"00000000"),
  8007 => std_logic_vector'(x"00000000"),
  8008 => std_logic_vector'(x"00000000"),
  8009 => std_logic_vector'(x"00000000"),
  8010 => std_logic_vector'(x"00000000"),
  8011 => std_logic_vector'(x"00000000"),
  8012 => std_logic_vector'(x"00000000"),
  8013 => std_logic_vector'(x"00000000"),
  8014 => std_logic_vector'(x"00000000"),
  8015 => std_logic_vector'(x"00000000"),
  8016 => std_logic_vector'(x"00000000"),
  8017 => std_logic_vector'(x"00000000"),
  8018 => std_logic_vector'(x"00000000"),
  8019 => std_logic_vector'(x"00000000"),
  8020 => std_logic_vector'(x"00000000"),
  8021 => std_logic_vector'(x"00000000"),
  8022 => std_logic_vector'(x"00000000"),
  8023 => std_logic_vector'(x"00000000"),
  8024 => std_logic_vector'(x"00000000"),
  8025 => std_logic_vector'(x"00000000"),
  8026 => std_logic_vector'(x"00000000"),
  8027 => std_logic_vector'(x"00000000"),
  8028 => std_logic_vector'(x"00000000"),
  8029 => std_logic_vector'(x"00000000"),
  8030 => std_logic_vector'(x"00000000"),
  8031 => std_logic_vector'(x"00000000"),
  8032 => std_logic_vector'(x"00000000"),
  8033 => std_logic_vector'(x"00000000"),
  8034 => std_logic_vector'(x"00000000"),
  8035 => std_logic_vector'(x"00000000"),
  8036 => std_logic_vector'(x"00000000"),
  8037 => std_logic_vector'(x"00000000"),
  8038 => std_logic_vector'(x"00000000"),
  8039 => std_logic_vector'(x"00000000"),
  8040 => std_logic_vector'(x"00000000"),
  8041 => std_logic_vector'(x"00000000"),
  8042 => std_logic_vector'(x"00000000"),
  8043 => std_logic_vector'(x"00000000"),
  8044 => std_logic_vector'(x"00000000"),
  8045 => std_logic_vector'(x"00000000"),
  8046 => std_logic_vector'(x"00000000"),
  8047 => std_logic_vector'(x"00000000"),
  8048 => std_logic_vector'(x"00000000"),
  8049 => std_logic_vector'(x"00000000"),
  8050 => std_logic_vector'(x"00000000"),
  8051 => std_logic_vector'(x"00000000"),
  8052 => std_logic_vector'(x"00000000"),
  8053 => std_logic_vector'(x"00000000"),
  8054 => std_logic_vector'(x"00000000"),
  8055 => std_logic_vector'(x"00000000"),
  8056 => std_logic_vector'(x"00000000"),
  8057 => std_logic_vector'(x"00000000"),
  8058 => std_logic_vector'(x"00000000"),
  8059 => std_logic_vector'(x"00000000"),
  8060 => std_logic_vector'(x"00000000"),
  8061 => std_logic_vector'(x"00000000"),
  8062 => std_logic_vector'(x"00000000"),
  8063 => std_logic_vector'(x"00000000"),
  8064 => std_logic_vector'(x"00000000"),
  8065 => std_logic_vector'(x"00000000"),
  8066 => std_logic_vector'(x"00000000"),
  8067 => std_logic_vector'(x"00000000"),
  8068 => std_logic_vector'(x"00000000"),
  8069 => std_logic_vector'(x"00000000"),
  8070 => std_logic_vector'(x"00000000"),
  8071 => std_logic_vector'(x"00000000"),
  8072 => std_logic_vector'(x"00000000"),
  8073 => std_logic_vector'(x"00000000"),
  8074 => std_logic_vector'(x"00000000"),
  8075 => std_logic_vector'(x"00000000"),
  8076 => std_logic_vector'(x"00000000"),
  8077 => std_logic_vector'(x"00000000"),
  8078 => std_logic_vector'(x"00000000"),
  8079 => std_logic_vector'(x"00000000"),
  8080 => std_logic_vector'(x"00000000"),
  8081 => std_logic_vector'(x"00000000"),
  8082 => std_logic_vector'(x"00000000"),
  8083 => std_logic_vector'(x"00000000"),
  8084 => std_logic_vector'(x"00000000"),
  8085 => std_logic_vector'(x"00000000"),
  8086 => std_logic_vector'(x"00000000"),
  8087 => std_logic_vector'(x"00000000"),
  8088 => std_logic_vector'(x"00000000"),
  8089 => std_logic_vector'(x"00000000"),
  8090 => std_logic_vector'(x"00000000"),
  8091 => std_logic_vector'(x"00000000"),
  8092 => std_logic_vector'(x"00000000"),
  8093 => std_logic_vector'(x"00000000"),
  8094 => std_logic_vector'(x"00000000"),
  8095 => std_logic_vector'(x"00000000"),
  8096 => std_logic_vector'(x"00000000"),
  8097 => std_logic_vector'(x"00000000"),
  8098 => std_logic_vector'(x"00000000"),
  8099 => std_logic_vector'(x"00000000"),
  8100 => std_logic_vector'(x"00000000"),
  8101 => std_logic_vector'(x"00000000"),
  8102 => std_logic_vector'(x"00000000"),
  8103 => std_logic_vector'(x"00000000"),
  8104 => std_logic_vector'(x"00000000"),
  8105 => std_logic_vector'(x"00000000"),
  8106 => std_logic_vector'(x"00000000"),
  8107 => std_logic_vector'(x"00000000"),
  8108 => std_logic_vector'(x"00000000"),
  8109 => std_logic_vector'(x"00000000"),
  8110 => std_logic_vector'(x"00000000"),
  8111 => std_logic_vector'(x"00000000"),
  8112 => std_logic_vector'(x"00000000"),
  8113 => std_logic_vector'(x"00000000"),
  8114 => std_logic_vector'(x"00000000"),
  8115 => std_logic_vector'(x"00000000"),
  8116 => std_logic_vector'(x"00000000"),
  8117 => std_logic_vector'(x"00000000"),
  8118 => std_logic_vector'(x"00000000"),
  8119 => std_logic_vector'(x"00000000"),
  8120 => std_logic_vector'(x"00000000"),
  8121 => std_logic_vector'(x"00000000"),
  8122 => std_logic_vector'(x"00000000"),
  8123 => std_logic_vector'(x"00000000"),
  8124 => std_logic_vector'(x"00000000"),
  8125 => std_logic_vector'(x"00000000"),
  8126 => std_logic_vector'(x"00000000"),
  8127 => std_logic_vector'(x"00000000"),
  8128 => std_logic_vector'(x"00000000"),
  8129 => std_logic_vector'(x"00000000"),
  8130 => std_logic_vector'(x"00000000"),
  8131 => std_logic_vector'(x"00000000"),
  8132 => std_logic_vector'(x"00000000"),
  8133 => std_logic_vector'(x"00000000"),
  8134 => std_logic_vector'(x"00000000"),
  8135 => std_logic_vector'(x"00000000"),
  8136 => std_logic_vector'(x"00000000"),
  8137 => std_logic_vector'(x"00000000"),
  8138 => std_logic_vector'(x"00000000"),
  8139 => std_logic_vector'(x"00000000"),
  8140 => std_logic_vector'(x"00000000"),
  8141 => std_logic_vector'(x"00000000"),
  8142 => std_logic_vector'(x"00000000"),
  8143 => std_logic_vector'(x"00000000"),
  8144 => std_logic_vector'(x"00000000"),
  8145 => std_logic_vector'(x"00000000"),
  8146 => std_logic_vector'(x"00000000"),
  8147 => std_logic_vector'(x"00000000"),
  8148 => std_logic_vector'(x"00000000"),
  8149 => std_logic_vector'(x"00000000"),
  8150 => std_logic_vector'(x"00000000"),
  8151 => std_logic_vector'(x"00000000"),
  8152 => std_logic_vector'(x"00000000"),
  8153 => std_logic_vector'(x"00000000"),
  8154 => std_logic_vector'(x"00000000"),
  8155 => std_logic_vector'(x"00000000"),
  8156 => std_logic_vector'(x"00000000"),
  8157 => std_logic_vector'(x"00000000"),
  8158 => std_logic_vector'(x"00000000"),
  8159 => std_logic_vector'(x"00000000"),
  8160 => std_logic_vector'(x"00000000"),
  8161 => std_logic_vector'(x"00000000"),
  8162 => std_logic_vector'(x"00000000"),
  8163 => std_logic_vector'(x"00000000"),
  8164 => std_logic_vector'(x"00000000"),
  8165 => std_logic_vector'(x"00000000"),
  8166 => std_logic_vector'(x"00000000"),
  8167 => std_logic_vector'(x"00000000"),
  8168 => std_logic_vector'(x"00000000"),
  8169 => std_logic_vector'(x"00000000"),
  8170 => std_logic_vector'(x"00000000"),
  8171 => std_logic_vector'(x"00000000"),
  8172 => std_logic_vector'(x"00000000"),
  8173 => std_logic_vector'(x"00000000"),
  8174 => std_logic_vector'(x"00000000"),
  8175 => std_logic_vector'(x"00000000"),
  8176 => std_logic_vector'(x"00000000"),
  8177 => std_logic_vector'(x"00000000"),
  8178 => std_logic_vector'(x"00000000"),
  8179 => std_logic_vector'(x"00000000"),
  8180 => std_logic_vector'(x"00000000"),
  8181 => std_logic_vector'(x"00000000"),
  8182 => std_logic_vector'(x"00000000"),
  8183 => std_logic_vector'(x"00000000"),
  8184 => std_logic_vector'(x"00000000"),
  8185 => std_logic_vector'(x"00000000"),
  8186 => std_logic_vector'(x"00000000"),
  8187 => std_logic_vector'(x"00000000"),
  8188 => std_logic_vector'(x"00000000"),
  8189 => std_logic_vector'(x"00000000"),
  8190 => std_logic_vector'(x"00000000"),
  8191 => std_logic_vector'(x"00000000"));
end package ram_prog;
